XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-(WW	_y5��}%�8�匓i-�����=fi���;���	����C��M�;'	��:^�|�;)7|�����Ҁ݀�kߴ�����]�1�#sv^HV��FmC!��QF(�R�q����g�(��ŵ���0���q����1	� �A�c  -ߥ�Qk.����Q��+�N��ȵ���	E(J���t����}�b
�+�G�ݩ�EOj�2iɿ�v���"@��Jd_K�UN=:�|�tXY����;�����I+E���F1����,^yOп�>%y��r:䷣7ȏ ���?]r��6h>����������-������r��΢�>�^],5
��3��U9aP>m�a�a�k�a&���Q�`۩�����#g�k�h�t@ϲ�AZ�K��?M0ʴB��T�T����yU���&�(jc������WZ�}x#B�z�����my[A�E�o�����Iy$&Ճמk��5��������n�b|���*Z�X��\,��Q ����D��C�
��@�>�����Ui>6&�hQ���7�}i%d^rPH�y��㡭�� i�Q�����st;]���[=�~DJ���(`�-ו��9zJ*>A�]e��x\�-ujKt/��5��8H�0#'������YL~�����@H-�����/:��3ML�B���*Y|���5���v��ޫ#�Ǝ>�!���-��O�&�E��@�#��C��Z�15Uq�^�9��(����XlxVHYEB    3290     c30j��ɢ����Xd|��\|P�����������@VJa��gf�u�4M/J`{�W�_i����15��})p��ݗ���F(�e)}-��t�K,�?�@_@�/D�,�9Ԏ�-ؑ�;t#-���-.O�MK�A�[��K^)�cA�������ӊ��}�sd��38�!vy�,`nQ�B�+|&���W�:�����������yF3�rX��� ��ޢܒ�`l�,U#B�[��U�Ō����0I�I�^k^�D�]�@�j���t��+i�I����⼅�	ΔqO5q4	mr��X���v��(�RO���e��ccU>�E��7�v���r�"�����B�t�>��E���,d��i]��5&��|��.�EeY����r�DT�w�����0�U~$P�܂��N�!qQ>�m��w�e����]q�=�c����|~U��V��ÃWr��JBT���Ijf;Wj8i9���<���S����=�*Z��x�����rDq�Q���l����Ϲ8�!D	�B�n_�X�үXJ.�X�N�e(���YΊ�;$�~5рZ�(d��e��S����j�׮�P�����t�:�ʄ�p�~��%�_�Ԋ����p:�AM�/��nV�A=pob@x� �Ի{�!z�J��`��:���;\���ߟ����W -	f���P�$^��l���|�l�1����ؒ�j��fO�.�Q;�[ju�_{.+;As��.g��܍�},e��4om�ù����_����ê߇�Әs���<��� ���Z�����k���*#�D�E'���<*�Ԃ�Aت���{)QXQ�,M�u�Q(�	pUؿ!����ż�}wJ����ؒM�^S�~Pݲ��6�&��M�������ĩ�f�c��;�{�$Ƌ�rש�|����7�����D�v�0|<Z�+$����7�M�-�w�����&��p���������Ϩ������Ei����Z� H��ȫ&"?^ ��_��>d��gc��^U�D͛���dCD�!�! 4�s�\kJ	]�I�A������Ǆ���b���
�t��I�I�S]X����r����1�܎�	,Zh�qݥg��lh�ޭ��1�V�@���������w]J�'
�!�L�� AqZE�SQ�%i4���v���a���	�����7]kmf�2��"schL���sU��0K�� )�\m��M��-��������h��"� ���-rM��
�u��M'�S��db�W�G�1��J��$.R�5+���L�;�����2�-B�:�ES��q@��Nx1��Eh�-K�8f����0�Z@7��JYT�Z �_��"ҥ}����6�2 �Un�5�:DYm�|�����a�c�Z~�Jr�Kj��\X�B�V(�9|FX4��Rl�a�N��-/�M��,��&[�U�E���5m��.%\�9�:�D��Βi(�?��S]�2��q�y�ZS������?�8�xWI��%��ِ�}�Ղ���2C��'�/��< �k�hS�URN1���N��}�P�B�r��p��F�^����T�ؿ�]\MJ�ٔVRYw.������|- ��fƤ����7_����C�����>��t�8��	`@�U���f�sJ��%�'}r���f�M��#�`�+�_�OS��h C��d+��g�NS���p%7�u	>A�<����b
��`�eױ�f�ٖw����\�[�
H#����V�0q�k�q���/�R���=��TIu����� P0ʜ�M�0�7����؁b��X��	Z�3L�1El�?31!�h�]�B�@w4���5=#l��^����r�D�p�	Nd{�uQ�y�LM&�+?��	�(���P�`8��,u���X��a�8=\�F��}^�&V�~�N'���I����H+/����M%�~E��xsA����v��6e*c�&�j�C��yg��KKH]!�9�p�m� �+x���QQ���X V�Hw��Ē�ML��a俟p��)� ���"�[7}�{=����,5���}� �"QZ�5��<-ꈡ6��)a	��Yy�܄K��{B@ҵ"��@�&�vާ���`�I��|ʩ��>�Jo�I��.���K-�X�7�)1I�_JK��)A�G�氩�k4�����b���T�~�Ҭ��g5{����D�.z�l�O�������(1;;��U4}�O�`u��q;�~ߚ���!�/[��-���(��P�KVm̛2� �N����Wo�n�z��#z���Ɇ���U�bQ��m�j��>�$Ѵ)�cF8���͛���߸��$�W�Ĉ}F�k4Q�a�:��q�U jX;��7(�&x�Γ)@��&���9c2����Z��w3�I�c�k���Zb�3�y��EfB�Y��̬��cF�-,��h_�7���(����@��d&b��?�&�(��z�p&��e~��u�o~�o=2loI�uy��;�F�������0�q���˽�&ݴ�H�l�J/��x�5��>�t ���5��׼h���'��d����]�5��Y�������ᢧ:�+LG�	����n��(�)t�p�,��H��ԛ�K����z�O��[a�U8D	����Te2���˗a��u�sQ	��>����n�^���xFP�kj#K�u�3T��pM�l�F�u����j9��p��5在���$���W�l���R���ζ�d��}����� M?���cnZ1~�0�Lm��D둶�P[#�"�牶S֣��2t����L�,2[k��Ř���I��$�7f��y�F@�JOP0���Ek�ԉ���6eF���66/�9qbE��Z�"#[�i�g]�XLv�K��Hɉ+�|�_�	c�W�8#���b/��?DqX� ��Ɩ$h����`b�}�ሉD��J���!���I��i*�i���DY��Y�e���N|���'�\`�m�q$��YJ�C�,O1�0���#���O�7z�L@���l�D���4�yA�>S%�f.P��	�$�mK�)���_�^�p�3f.��"<�q�