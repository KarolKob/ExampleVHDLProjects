XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Zi52va�.)�R(����UX"��m�o�r������1�t��V5��!#��v[O�����z���Bs
�A�VJ/f��W�@���YA�Pn��X�Ѧ���jh0T�	r���*�����O&��0�$�]!�9s1z-@�����o�6�Iߠ��z��\�x�=:��5�gGe�5VśjE��x�?�(�w�������-m+W? '�*�H��v�+�V;*�}��٠��=�j������8�zP��l�Q�[�O����j�#a�LI���x�Y�G޺���ʘ�8�y4l����T�7K��Nd�;�r�@=�؊��8Q��%鮞���u༓����.��+�~1Y�*�=��{ve�p4�P�}No�"�~p^�X=[{��?���W2��9�����'.�k�i�*\�P<����!�;Թ��XF�S�V&�Qi�hQrc�7��뎋��M�˲�J���08�h��I襁�g���G!#`�s1eE���c:x�����NL���Z*~�0����l��**	w�"�ԥ& �u��2�=�vn?���E�|���j�wߜ��<q��1�K������o���&�V}�w�&�=A���0=
����x}D��1�Йgc�mC�T�]���D"L���V�|"�D�kڤ#�?��vq�����)��,}�q.x����9���
�6ެ7��x�W֬�S#Oτ
e_�[i�a Ġ�@j�N�jBɫ%��U�Z��2h��6�#��XlxVHYEB    fa00    19d0T1^*^B˄n5�d�zz�h�����d<~UD���9t��7Ε�k`�󐦔�(��Ju���g�b�w���,h
�����h|8��aB:8�g���&�A5_=�L��Pu�) <F��분���&n6�Q�4DKJ��EޭS�L�h��r �� ��H��ctٖ�pޜ��0(E�+d�6�����'V�)V�f�|ؓ&"�w���CZ��O!yP���qx�N�3D�ˋX�U��uB��.Q4�HJ�ó{�I00�B������:��BW�6�J�E%C�R�G�b(�9З��ԭ���I�!Ȫ7R/�8e�t��������P
��L�8R1V?}�&<��p;O��9��i��
��B�P��
���,���ī��x� �Zd��@�U���5:'� ��{,%�:Q�V0�w~�F�*#XК��D֡�WM��Zc��0$��s-�)�B�qkI�'�l��@�f�n�}�4�f>ё���Df4(8�ޘ��K\pB�h���0�!�3����l��`W�]uI_s`�R���|n��R�(���Do���^a���3R���� �̰0�����9o�&6�V9�R��ʷc`Fz�Ŷ������![eH��������qh�K��d������G�*r �wD�
�P��0)���b0d� %�ժ〲�������c	��1�VP7�#�뛳R�T�W�P���F��Q����GU*�Đ��Wj �"�{[P���GBS��M�8���t�)�%f���[CY�T�s� �{����H������S2��5Ķ�M*�l'�~���C�Q1Hw_��Z-Й� ��~�񊔤Vu쯱`v���aYm&<G������ȧ���3JΒ)_~�2�@-����7�^�/�8�Qѓ\cv��;�g Ӫkr�$J�(���L�6�Eٍ��_�X�'[z��|���٥H/��Vb�q(X���6 b�R�Pi�2��{�,�߄�d�A�(��=t5҅���Q@��[}���3Ҙ۝?���6��ܦɇ��.��x�$)l�g",R�f;�)��fG�n(xF��.�!���kd�m���T��%Q���m�q�r9]ILl�����S ��S�ǅ2OM�R��S01��v�k�y������2���z��	N�z������%ʻ���C�/�L�,�([]f&�ç:�[�25� ԑ���0�W]�<z�t�Y/X���|�0��u�M���o}�kf5�_9���h2����W[wd��i.�Q��/W�P�B�l��2��9��W�}�&+�Pl#,��"˨Ĝ[SӸ瀀sm=Ĩ^8M;l�Gz ��yC��t4�vH�G�A���B��Q�;�}�3���
=���̿��L�yHpP�x�勦A�?�+s��7�U�_���R>����(Y �zO���0�Z��i�+�:B����6��ݿ?�c �Pګ.J��w���&Fr7��?V�spE��mӀ\�Y�V\+d��+��hyn�u��wWC������{7��<!X����^`���ߟз2*�߰z�~+��1����DZ�tQd�	�1[?7vj:/@j'����R�d�a��,jv/��Gk�����~1;�{���Y��y���༥��C��M6�����@25�g����'&�Lρ��:�͍�Ɠ��/���5A��G����`�s}�p|KA,�(�n��{�>�a2���� �/χYK$���mj��S���S�Y��p�2��0d��L��B�N}�j���L����4&]�L
/�'i�o���)&��Y?Ԋ��R!�(z� $Ř:T�x�8c�Ih4
�R��_�$@��5�FN�2]��z��ZK{۳��}\n8s�ױ�T�!k=�f�{��W�j�ݾ8K4����'tB���k�kЪ���>��F.�ѽd���o��嘯 g]	M���&%RA�]ZM�8+��,(&��I�O?GiV!���͎JC�B8�]N|Q��h�YiI_�ƿ­�q�$��w)�f��~N���O3����ء"$,T�ݸsV���ڷE�會�4+o�Bƿv�.0�x�S��bm�R��`F��}7���ݳL4W�����XH��r sp*\��𬬚�1���� �O4^҆P��ҍD]���-��)�<X��&���;�2I;8%�����ſהX��Px�n��A�O�Q����A�����B&/s�Tmo z�km{6���l�n�O�Ku&�����^/_,7�Ѹ��<��[�9qwF*�D5�]��lO?:z`�&�QO,��Y� �T
_����xYYu���fj�����R/HO(��38�	#<ra%�
��E��I-�7l�� ����Z�l�}�ŪH�|)�:�r��꾟Yʂ��"�8��S݌�q���3��ֿp:���ܣ�&��x� �Ѫ �L�n(�p��n�����*:lF\��Xd�j��Ma|������)ے�0���ц��V���oC$ș\.b����k�K3�^��^S��#�4����tFK{?jE"n}6��ƒ�U�C~�{g~/K�/�6i�(E�:mT{��lw�y��k���Ѡͮ�J�^ӯuR122���X�P��������Wa��FD�=��_�/ s.�M�n��s�:i���&|�HF�� *�5a]��������B�R���"�U����߻�ǍJ��H��^V���m[�D���f�����M=���S�xNŐ��j�vt�4i��RD�mY�I��7�!6��(!(�Do���8�=e[�2h%��#�WG3&.K1��e	�@����__�ȍ�8�0��&��p�Z���?��/�d{��sh��7�v"&�{#����Sxat�ײ��d��8;t�A��\*ҟ��걉�G���W������<Owf܍��j�d�����S��
�����x���̤�����;��&��m���\���wh��^OڭWq��/��|� ��Q�y �U�3��ZSq޷��(&6�#�x�h�Q��b\ޠ̴y�:����~�ilz�`WΞ�Yr��X?�� �ULÃ���ˮ9W��"�Qw��7"}G��6��þ��A�.��2��^��I���/�G�d�2��v&#`�����ڄ]�!�~��iQ�&���&x�� 1�.O�I9
���v�r����G���i��?�s�����5�/>u�x�Bd�o���ͯM���C�|[��$U��!0�wX�H�ODc�{�z"�}=��*�@_������ۂ,�b/��!���	�1V<dA �>`����U�=Z�xV�]������7L{u+t�X��,f�y��R�W��g���Y�c�Bf`����6p}�;� ̒�J;&�!4�>�邉A�כ��.����Qg��Վ�V�kv91@��?p��K�f�N�Q$���j�M�N��E�I�ѷn�B@0Y����>�dR�OƲ)�F��?(��a��Yj�i����\'����E�����x��#��%k���S{��l�Sa�o�H�lJ�Fj8�_��Q����"�9��M�ʣ�����k��Ӄk��H&[�mX��9�\�QJ����*ʻ������-�uëROM¸,�@��!�<
y_��)�܈,2\����6��dY\�Z�&��Z����n��%}~AH4�P�O>��k�B*�ֻر9K�����s������o`���o���_D-H*����dx�p`�0[>����A�-6�y��q��^�]V��v	�:[�e����"�*�2��<]�C^�,�\j� ُM|p��u�D˭�l@���`V7n. �*��|rv���ê.��qxʷ�^"�,�t���%RP�
��t�[3��F�`H��EE�
�C��k*��� �]~j�n�FFBΥ��=+�og���a�1ˁ��7�����}]U�f:��K0�t��,=��(.����|�^�6�������1ѡ�#v�3���$��
x��!��C���a��+��UR8ܿ2rr�oI��̈2����{O��A��~�G�(8��������d��42і��j!�G�h_a�dD3���m��J!�.O0�� �����s���`q�]�ꅴ�����S��N-����.�������%�y���-D˟��s�|<O��;�^S8e���;���b �N�D����4�܏�W�I^�Lz�-=C<�Eꍟ�D��|@����N�*���y-��e|I�#z�#��M��	�F��ջ'��xN��_���:�
��=��Cq�ZƵ�8k�t�<%P��Q�V��us5����Rʵo7�,����k�����fwۭ�&�������7�M��\�,����E�Fm�3�lt��J�Pv�s1^���Lp�a������<eG4 ���j��:��t��{f��l���&%�&�����RM	
�A���'f#:\�iz����aek���V��8����'=2Q.���o�����#�ȺZ��P�U�6�@kQOM"'�K���$��~��h*�����O��!Bi���L5�~E���	(�$��W�C��̊v||<�'���[,�!��tPa�ڃ^�*Hfn�ˉ �d��L�:�ۣP������A�y"'�Sp��ʵ��)٬�IрNo���b��%SVL�Y�E٤��'���^�t�S������f�'"�)�vI�a�,��F���p)!5���F���J��5E���>�]����Y��*9��Xܿx��i��V�?���7�L���u�U#XH4`}�G�����jc�1�����w^��L��E�rܮf]�<��jX�W�a5(�Nxꌘ�Ι[�4�v����cZ�Uy�̨����I+6F�H��p�岟����@�-�����Y��m�@�H�*5���L����]{�ܑ?����,w�,�a 1���І`18���L������ZN���hc��փ 3�SU����A�F�j���/�T>[oj�C aӧ���ַ(@�ޞ�.�s�_;��}�;d�UWb�9�������u�*�7�����-{D��d���b//���U���%�A�=m4y�fr�8X�A
ͩ2?� J�>�}�i1�?F[D�nE�����a�4����?�߱k}�M�t�&�OI^��M�~7㛅nD��J�[wj���������b�t�c�c�3��j�������®�T�tb
��[�o~�w [ܞ�#x��||?GJn�X�:E1/Q�q��c?�����(@� ��l�D9{%�ɜ]�qpr��n�' ��H(.�v~����?||8��6	��1�9���k[b�0G��>!#{|��=���]�Dڔ���!��G�ﵵ;�?�	F�fc��=J���l@<���-
�5�-�3�m�#�9Yi�r��._v�pnY�j4��v�����M��^��Yλ5(V[��Ќ��.TnWp��� u.�
P��4*�����^��wDٙ:T�(��g�hx�L9C�W�*pj�X�D�v�;����n��c���)5���׵����L���M�ș�X��}= d�7�_5��h���������k�7�P)�,���?̼�����C��U��g�.�=QKZ��nl�Y��,���|����Q��n!��}�xH�%�{�=t#�ٲ`[.V[���%N�Y��G*��9�3��n��4I�Ȕ��z�����
H��;�Zv-�$�uɇ�T����%8�19x�Ԑ���t:M��u'lG����S<P�H��DF=��{��"R� ^�"����H�?O�X`��D �ݮ�������;3�Jw����B�ou��B�l�L�b��5�� ��G�����'��^�1���z�Cw�I�,l=�Z��7�7W#���>D�s^� LP�)2E��{����7�:Pm������I�!u�՞��-����H�������]�ap��"
�XS��ajq���MQ .]@��ț���Z?�f�ϼo�m�8'}��a�3Q��W3����q^�b�T�Z�D�^��=f[���E�cS�R2a=��p
 k�A���J�R`�A4n�%����G��+v���	$�m�Z��4^�E[�鄮f[a�'eMA^�ٓ�	W&���/�V���,*\YG�jP��L8,��-��f����I����ya�^�>�L//����_A�n6��ڏן��#q��F%Rw}G~�����Qh��@%��x�(%_QVL��B����h:�������Ny�r���Mys���pG7[Z�F��Y0��?��Ϋ:u��C�� �۰���r�7�(|u�VS���c��	`�.�P��1� �B����w��MH�cy("
#��(���H��KG:�d�Z����b�<)+�%j?����~���.b�w����Z��5!DD�Srb҂W\~Z�:ZJ۴(�z�/� ;�V؍���o̷��πp�c��ė��y"���\�,� ��.�!��,��2�\����&K������(Z櫡��fv���쥃؞�����v�6rXlxVHYEB    fa00    1630&�䁲MAW�uܳ@��qe��A�6u�-�}�;�¤U�N|���##�H�X;�tTr�������Q.�G=㈏te�� YO��|3�gՏ�@ܥ]��h���e�J��H��p�%�9,R��Ls^�r;�ME��6�>�du}q�MLS������lj^�ڡCm���8K�@�����|�h�1&l7 ���L���� ( �쌚T����ȴ���7� �,�����̍�������N��J�d���uuv�j��֒Ķ�[�/��zŢ�������G:L�zd�j�'���;7���Ɔ��u�2�C�	#l�8sU����E�W%=��彥�w:��8@��լ-����_�#�;;x����Kc<� ��e�Z��o����؜+�%h>�_ T��ǰd�ԥ7�j���^IF��=B-"fQ���KQl�.z�qZ[4Q��z%�Y?$TAF$v�Ϸ�̄8���D'1�Dc�B����U\5��kQq*�*���@�"������E�~�,���^��!�^n��L���}���諫	�q�z�5��!�ǋh�Ņ�EO����`i{��?:����Ӹȥ�)`4C:E�DD�����0�
��t7XReg�:nC���Ͳ�y�}�T`���H:?9�K��ܜq;�x_�&eHJ��}Ȍr�V"���.y�&%w+3Ap�m(oz����}����ӕ0^MG9㼑JJ1�i�����G?@�Afdt���Ae�%�m�
��щ�_a�a��/<IH/�i��>�:�~��T�
���`}rJ!��Ay�Gg3�oΓϡ��v�S!̹1���Յ_��m�&:䵍���k�
mJ�-$��u�V��iO-�'�TRg�v���<��̌��"M�@8w쵑pu�T5��{�aI���/�Fj<�h�j7bH�~�>�]�r��8?�h��RJ�:�A�	��Bd���>?��yA�i�K�"�����������ܨ[[̇�+�Xf����"}�Tw��k�(W'w�tOO�M`"Ą��9_P=�=#�����ۨ��K-Z�i6�\���<E��n�ʸ�짅�N�S�?/~�^-��S]����0��~�)�ռ�X�*)���_��H|�����!&�B� ���r�3̯�[TC>oy�`˾�����z�г\Pi�H�H�kJܛAP&�G��#�|^i���l;\�Â8b(�Q�׉^�g\R�Ԍ�9"¦n�W%1f=\��x9\��ջU��2�-"1a����\�ג�}�Y�E^�iZ$�>���+��&VM�<��=���:�T����ݧ̵$�Xc���1�
�y�As�|6S��z���	U콭������l~r� �ǄO
�H0x�MZ�%���,�H�ژ�̪����9���Gp_�(sG=�I)��ˤ�R	�d�� �.��Uu	��>]��Nv�ǩUX����]Jn{����1���tL��}���$�#�ve氫�x9C����V�6V2%���|^��9Ժ&5]�r�M�e��V����s����K3�C&2	j�0h�T ���iT!t7���f��k�`1��")��D�Q����CU�"*��Ec�����3��<�	�4�aM��l(V���#���������I��a�b�/�O�����0A& f�	S�Vu���r&�a9��=��Y�'cZ���b#Y��n�n��:{�������?E�b��AG?�x�笸�׏'�u���C���_�qӎ*�F��A:n�a��ۨ:)g&|�ɗ��}nQ�	�÷��y��/qo[�B��?�_�9�z)��$/bz���G��<�v��^�9+���y�|��$;:U��3��',iG#�l���0FO���O2`(���[��z�&XN��h��� ]�6
7�����A����p��Gː�!1#aj:�tb5�����	�Bc��v������r�q��cVKv���9��yP�<�j�/��<#=@�;���J�Z�W��+���o��T�z5�9!$���l�D��^��߳bD��'@W��A�S�'.M�wfe8�Z���"���G�l8.W�snϐ�U��m�Q�7W0��k�
Fqe�W`�ddЫ�)�z����	��q�Y���e��A�n�m;M�N\�Ψ��(�K��( Sa��9m߃��*~Ä��t�zP��m��f��rL�����3�a���d�E�����fDbL������5����LL���ꎺV(݃bm�s8�e����s��|��7/˂���6P�����zg�5���PFp��=;�K�?Rv� P"UEM�u�˔e"^=sU�:�����\�,��Q+�]�i�� e`v`�������Va�RR.��f��G�T �-nU6˖8�Χ]���^�t��P>晢�b�g�����c��څ��Qv��a�"aZP�ڑ9?�����6AS�Ii7�뇥��x�9?Z�RGh�UQɖ8��q4��mE:ş�#�#�y�K>��@&.)J����<���ݲ�f��Ɩ��_�L��ךּ���.4�Ou@�w��=͕�{�ۭߓ/V��,^#U�%bͶ�����Ww]!7̮^���퇎5�֚	�K'��pf��Ve���/蛺���@ޠ�zꋃ��7�q7b�������>�Y����q����+)"���1��Y֝8<�ay��D9��X4aC8�F�	�7$2iαT���~)zOJy�8Ү�?:�O��Ε�ֺ���ʩ���=��݌%����g_	&L����2EG���1�#��^�����`��&{n�0+?'�mZU��ނ�C�Hm��Ӷ}$3��%����6*��ë�p����iiOU�kɔ�2���İ�@W(!�1ο^��K�[�U7�]P��;������xI��G`&"��؟��d�����S�Ī;\��7+�v��}Z��^�'��PQxL��r��L��#o��I9��d���=����d����N�j5�΢����UwR[Ɠ,�Z�YD�-u_#f-3�Űh;�[{�VfF7:C��f|.8���*R{z�y�5���#� ���GtS�+ߐ��͢z.�9�f
3g���K��apJ�Pޕ����P^�z�|i9�S���7�0��W�b\�j,'���G��i�Fӄ��Gر�ӈ-N�AB�����^�����d�t���� �jA	:�q&����c<_Y��D�����3.
�8�ֹ����i^�t��QH���С������L�"pesw���x{���SST��b��?�� @h�h�ⷯj[zU�&s��
G�Y~cG3H�@f������|c��	8]�i1��q�����d���D����>6R��*^���<Zy_VBgm�-��O<�y��b��������=l2�O���Q�d�T����E�b;o�ed�KpI�FNF�=&���ef"��t�+�Ã��ih1Yə�a��+\�i��C�d����A��Ĉ����E����Fb}[$����y��wAO���c�<ų�i���Ϛ �N���Bڕy�<�Ȍ��p56�ҭ�ݾ����&��ӊ[��]A+�#z���5fq'e��v2j"�]η�?"v��j��hQ�� �3r���覩c��f\�I�}0��|���\�Aᅹ���`a�ib\
�}����.�J_w<��e��[g�RF���[������{G*�!"��=c64�	3:�]�W\����p��B��f��TA�d�5���]M���h�	F�g���`�ǰ�fV�A����H��A�k�B	7��&ݶ]i���%Xٓ�u���{!�p@�a���v��`&�9�_�j
���ğ"�U�`�6j�r���C�ʖ������{Ɲ�4��q���0t����SS����U�Z_C�����G�$�=rhs�t�KS��,r��9(Gn�8~�k�g�4�zG��G���^�T�� ����}x��D2�8��U��,C��1�P�Κ?t�Sٱx���%�nq}�.�S���X�$�&�#}ڠP�
k����=6�9�J?ܞ��䉑�#�IQ�e{�H���?��_C���QX��x�"�t��Mk��R9H. KzO��7�)��+{�h���CAr�X����*dj��qd��}�Z:�W���MV�V;ƹ��U�u�f}�&
t�E<�r�^����l��
b�;��#d�ڢ�{�h�,$�����u������Ɉ�����|9XA�F֛�:�]��ޅ4&�?��;!T�;<Y����EV��~��/��`F(e�~;��4�q�V���*�8�IE�9.�� ,��5�k�瀚Jq$I��.7=�vX�^9�IW7�U���5k\g���U���b��zW�����[޾��b�K���o���A����Eti���{�9�������6ʗӴ���oG��x 0����5]�����y��i��B�_pLb�tU|�P*�ѵt*O��(H���op!7d-lڌP��3&�d�a���}ZϿ��<��,Dz�}]ge]���~i@t��n��g^���/H�m����%������v�L6$� pt#T(���ܾ
~hd0e������[$��Ml(�W<?]��!s��k�\�F���<�����yY-�����2�;,���7e�
���_*P#"
 z25/��5���"�6Ϳ��ޚ4Zɨ`��X�Ǘ�!�$%A�9�����$��v��y���q�*��1�K�1}�T1F�]$���6�G�ØU�x�s��>S*�kmGgݜ%Ubn�?������/�����"�6?L��rPr�L _H����پ�o���;���[��ʍ8��*te\I�&���O�9���|P��,^ο�-�B1�4�״���.9�m3����y�mw�\,���$^6ŧ�<��He��0Z�����T����Uze�����W���C*�fn:]HWe�.�'�qp�[t��UJ���H�3���<�:~�����P���Q�].�����u7�a� pvlK������NDg��c��sYnf�6�4Y~\�ɭ����ȂA�N	��I7���Z��ԽV���k��#kl������D:`N�m,�u[v� �sxwڻ�;����"�_�~E�Mr�!�1���05�O�`�#��9�9I#(|^��{���%�S\�3$ߣKs�Ǝ����;� 1A�b��#�?�� f)��H�Z�9�7 �`SPR")�;��f;Y�`�b"�U����U-��gU,�1Mk�wd��1��'�Nς�+A�`��o#y��9H��C�@50�	o�'!4��@~��i�;��NXg��)#��t�h�smtFv8��!�Q��l��`ge��I|��<���lM��W)Y���v:4aS	5�@)G��0��36��e�[poh�O8 P�����J(J����{�[�����*幤,q�c�_d����Y:c��~Ր�vD���R�%;
����� �@��n�����ک��q����S'�^���87wY��Z��U��������.�i�� �j\Y���Xr��XlxVHYEB    fa00    16a0��K�i+�^���K$}K�{?�#�A���hF뱍2��e~�V�Cs��DG�?4|�n뷵���a	<��L��y:A�b�F�� �����EaA��C�ى�;��2�g{���P��ܩ��#\^Y��ګǗ`�@�b��^>u�������W=�vŮ0�5�Ng�h�@�0�'Lj�a)6���{�y��(m/D8�J�w�����Ux�{E����}�XZs�C(�iD�ru�W� �
_ ���I���
���YYϗ��M3w�3��l�\BS_�:����w����x����(A�fXP���UY,k|����tL�<�vGa�!���[[]4b�DP�+z�,VF�|@��Ei�Ó�@n٩�e����Vx7y���ַ���� ���V$����1�*kmL�{��|
|��-�T=�ԩ�Qm��Mo�� �_���#��٫�Z�p��H�
@#��g�k���Y�fThO��s8S���aOW&/�	, �r� F ���'{��/v���T/ i���޴#�=qF�o�&���I��k67�<��=�[�.J�c���h!q;�%w�V/��O텾�2�_��"�Ǒ�tcnK����\��{��M�[�5�I�DECOjc!z�����m�	���QM���{N�{ʴ]�3b�'����7C�x^��^��>�[��Y�wk��L��5����X�h���k��C1���'�G�AQ����B��n�������F���IǺ�4�U�1S�mj��&�b�҉JBujW.GLF����\r��4~��#;�1::�|ƶcN�@̽�����W-t5��TJlD�;�?�n1�͝`C�@��AYȔf��`�4O��1t_�,�U��@U����.|28������:��഑��n�Si�3��o.e(�(��Gq���
�w��y�t@VGQw:�����������}��C�wV�u����ä�.��D�qX�l���-Z����U��q��F���b��R����UH@��q% ����{P��*� ���(�a�ł�^L؁��e�6�?�����}�%�j��sS�!���-�v����oB�Ki�pF�pQ�X��P�Zy��7�R2�.����i��r���� �/d�X[���i{ϴ<��
ɨx�dP1�ݿ|]��r8��q�Ki����sj̖��6#�6�_��E�)z��G��`�Jqw�S�y
���$���"��\�ȇg�"N|(-a�y@����H�b�����pE����k�ob�ɜ	܇ޢg���R�l�}n֫�5ia�V��sb��ݻ�a�L�����a[��zĕ% f�m?*�-~�ӳ�݊jC���GV}.x��h��k&��[�W����B�d�2�E䗩1�������0g�}E!�\X� ��I8rt@�g1�+�t&&�N2���L�!�7, ��z�0wl�7�K�gX��)åe�>�J��Jc�����Ju�wGuIx/W��j,s
\A}(���D�� G^eo 	���:�;�)ه���i
�piNbM�)��53�D�k���,K)o ��_�7O����o�g�P˶ WA+}R��)����uFZ|�v[]n�0�.��Y_O��a�P?) ��,�/��vC�!��zW=ʯ�9U�\/O�M2G�l��j�1�D�ŰON T�D�����*�t��v��;�Up��z+V��*Qu�+>����MX8$0�BM����w݄��lT� �#Lp�م�M
�����	W���T�Y䃴�k ��� �!��ӈ���ގ�|
	z ���+�QY����`B!,�X�܎�9�G�
��]�(���=	>��w�|�~Y3S	Z��a����Lh�O.�L��(���;���R�k>��S����&�#��×��X Ț�M����!{=��VU��āJ�0�:i_����l������Ѭ��*1e0>��A
<������l���Pl�j�����8�,��j�	�sO��J�[���I {�b���C�߳f݄,8�Px,bepC���S%ռ�5=RZ��- ��Eg'+Nʂ�0����qf�p,z� Ur��� �N��=D�z��K�c�>��,��]ҁT''ƕP&�i}u���m��}�=�m�D��S�0�CZ@�]3/�q����;�ko��<bm(ϲ���^:Cg[`��p���e�eb�eL����u��߀�K���Z�ϽIY�ko>�Q!~��r��b�+(3�Iu�=�q2A�u�Ur�����kk�����R�&��8�h�d�ݖ�<�D����ԩ��u*�n{3�?[�@N�Wɤ���rr�2�ן\H�B���G�f����p�A�Âd��.`Ӷ��U0�,��pB�c�$t����5e�@��Z���ɭs�F;)�r�co��U�o��4�|<��4�N	�ؘ,�(���d7?m��ӆ!�������Ư��W��x)'�Ow��7&	8AM��f����#���EW�����Uc�@�,�<�*D�Bgd{�OO��@�/��i��Z[�D؀���'o���֡�ѩ%k��jh�%��[��n�@��&}tblR�5�f�߯A�c%>�.6�I���2 �$����-n��wY�&7J���"�_�EKG"�G��-4E��s����c)�"w���ᄅ��̟��l�����5%}I��r��E�ȶ��O�?x6:W6a���J^g^�̰�� �i��OA@���O"iC�u"�cdK*�t�P"��4l��#"�K�+ZJ��uxf���N�"�����_��r�4�ַ��l-b��x��r�F��+.�����̄b#�yvv��rPgyA�_�L%Z�@���O�w��>�k\,B(����1���r`g�I��S�^"��m��q�z泐u� ^�����e(�n���m�((�)_�A>S��+4��EA���9+�tډ���u'�H �B�O�@	i˦B��Mk�^�r�������)�L�x����Q�o1�p o��vpK71`(nL^ꣶKb�QAs�M�kU%�����ZvS����ybAX�����&�EB/�}��#�U�y�O]v��!���(�'���S�n�42�'7P��ǏH�AX+�����j̙��� N<�Л����o���|�$���qRAh�f��^���h��)�k�
��)�|�1���s-��Ref�:�2�Bc~ے��ʢ-������NϷ�L[���p�Q�Z�Cc$�xA��
P&�3��gl�d8lP �^��~8ɷƖ�\� 3�ۢ�yB�ө�� Z�zw����1�I��b����?��B����#'�2�2�����Q!0��z	�u&���m�ä(H��9kHf�5��T�X�:�@ ?�]��/�lSPuX��_�u�A ����>��"m(����X����`���8ƑO(�b��1�=�oWW�ɽ�Q��G���7�$d��g��.b�?"���Ey*�2��k==�����#�4�˘������O7�f����>�0�%C�dC��)J����F�ȗ��	�]�q7��������"tIn�7��J������ڭ��z�pU��k��ł��t0�y��_U���N;>��^�_dɳ�y��+_��������}~q�N�R�m�D	��0U����q�#��� OXZz��^��'�O�a���$���<�S�[x7mE��ĲQ���3�#
;1-n�����LTԀdX�M��y��#:;��t��3���op��W��\��ˮ��K�#X�"�3r��;�yK|G��H4O"���5	��̊����oDtsH�)Ǝ���|����2k�ܙ��O�@n�!TK2!��n9��!���G�sh{"?fp��x���K�f��� �Ԕ���Y�������-�?������ Q����B��tȷ I� �e��Y5�:~1�m)���e�fʝ��d����<�7m吖�ٛՋ��0h'?:�z1����#��� �`�����Gf���L��Ѝw� ��E�e e8�������Q�`��^�n9q �47j��X�|�;�${P���;+�8\� �`_d�/�B�� �L�$3rj�3I:��R\����|.���r�.�5���8���-¡os���[Ё�q�s~�<�U�j�<�)V�;���6 )\͡[��uq/p�E�+(@5��܄(����țA�}R��aQt�hI ��Z�~���Ã��}��ގTf!���K�Y��H����y��صLY�y��}}��mg����2��ٗ4�v�P3�ѵ�È�zI:����_�!*?K��p��W9�<ei���L�5��u��Z#��<.]����x���"�6/m�r�"v�ɡ���x�d6��{�i��4��>���+���pޚ��8����#[������:����AP`�?Fs����DS�'��S?[6�&��="$ht���]�s���Gw��Dh}��e�Px@�(R���aB��1��=��S]����T!|�� ���8j�ą�`�iޖ�q=���J���D�#��i.ȎZ�f?oCe�,1a�
;{@�MO�����ʪ�\0�
Rv.�=q�u9����^�	B�ɚ�@Z���4~��\5�)r���5CS��T斵6��E�@q�㥋�=�EA4�5��"�+) ��4j��J��k��N�;��Js.�T-���yly꒰��3�Giʐ1��_�o��m�_u�+=���Y�C���5>R[[dc�?<������{�Wr&����޷�^��Y����>B',�7QA���h��6��P�R?��W�ۈ��N�8�[B�y���%�̑}Ty����PI�tU�,6�JY׹l"��%�w�I���I���./�~���W�/ަʿ��.��D19]�}��y� R1��	����q���
�q$���Uk� ��%��/��qy���v���G
!%! �
 2����k�	w�}FLh�m�u�R�o��nGѭ9� R-O`~MJ����bj���Z�}�a�}�5��rgi��L�����ȟ��|��i�g��~�	���r${��A����-�����V[���ll-� ������*����B��(�KT�p�F�@os��X�M��2��w��d��W�&3 ܱ�=/\���8����$�������	0}�73���.[�������'�� ��_i�0���b���.Ҫ!��XŴ�<��%��~3;�鿡+_��ݠ9Pq;Q�����.�=�k7�x�K&���̑��&��(�Gu��U�Y���K��5{��t����b=��,.����tv�j'�&��|�՟���h}�Z!�1Y�c>�ol��j�b��X��|�B[�35J��յF2)�����
�v�'P{B�[�N��^�zk��B���W��>��WG0����M��m5&")���X9z���J߭AuIL���n���a+�W]T(�.����IV�*;��� ��mO0�l�"etZ����͙D�n+8~���o�T��
��Iݠ�GR��0c��a��C!�g��
"T���F�zᵠ8�2m�n�+1`�ь��Ұ�������č���0��v�hjp���FR^<X��K(2#�%2i��U׬���Z2w(XlxVHYEB    2889     400���B�����4�C�j9��5V������T���7��^���+���7�cƩnb)�R(D��`娄_h�8�M!�>{� yr��p����:s�͌M]��Cw_����
7� 4<A'��U"��z���*Zj��]D�����B7�?=�N�G���7��}�����Z/��U�8�"nsf��I��v����ycX$��e��k�����໤c�F ��^�)�����m�r\�'�')z�Ź�N�_��~3�(2�(��;�-��-I�|e �|.�.���+:8��F���Q��U%�C���7�%�V��*Ag\�$�jΛ�J�"tnU��	H%��P7�K]�Y6q0��7#�Db{���u	X�]aT��=Ҥ�T��^t�4��>�u�V�C3	�ԍ����;~������ڭH9	2-��+*���jo�$a�E`����/{������`��x�1�%�3�A3lh4�����4�RI84 �G�&����]f���RFǖ��H&l��0CP��RSd��I�yl\n����ttg������[�;Gw���g������t�X(E$����'̈́���p�XcS�m���[���}]8T��+Ĳʊ�Չa׆��>�J(K�.���6-SYF4V6m>���dC׾�r~!_Ȝʇ\��T�'7ۑ�r���E7è�p�MǙ��G�V���s���V�L< TD$�l�Y���$e7i��u����������� ӫ�r�"�N:;+�#d6�>q�	:�ڟ!DLq�-���ɱ�,>͝>s�x�:y9���]c��n���l )��ā���gqu`�"80��O#D[͆�?p�o�D��z���3��/����kg4��=��/�~4�W©lY������VR�kd��Ǫ���I�d9'�)�q.�+����� 9�eZ�$�_��4|���Z�@�����8��H�� �WRK��Yw������o�q�  ���R��$����N��5W�H~A���]�C�