XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ղ����^���#�On�0��1�_rǵ�٘�	!W�p�8�����ʓy�n���jx��?Ȁ���c�i{�E�b�#���!x��?c�0��2b�T;��j��wyQ��7*,������QeDH�j�#u�)����>����r:T�gmy,M�S�gcf��a��UV��f/ɶd����3M����Y�~�W;N��i�%م��$e	A���2R�\�@��˨��� �p�s��c��Ig��y͙O�T������#%��y�֤�v��g_L�S)�
���w~���.��9}��ºi>�O^.�Z�����m�����_y��eο��-�+D��RE��#\G������ �ǥ�Z�8\����!�4����X�5���n�*����aܽ���������.�����a�Y����f['�K�.��B����*2����)��^�w��I�X���C��&p*7ܽS�@�	"'ENϖc���2�@�XM+ʐ�L�~Zb�S=|�O�Ꭳ��%
%S*XX�`�&*Ћ�t&�nY�*M�����1{�|�����L�8�r����< ��X{���rq�eD� ����<wf�>�U
�Z��}�r/$Ww�)y�ְf�y��$�T�1�:\���������?;��iJ҈�p�{ ֔��4�AG'���>�9/��=`4xy�.&��t��7�q�by��ԭ��oɐ=M�xHvW�~����}b���z&�WR����H����u%�H0������_+���XlxVHYEB     b2d     3c0L��C��{?R�°��D_�G;�ވ�^����(�[��"!{�{������av��2W��Ձ�ٯ(�����KgzP��iI��{~�ܙhȽsZ�$c���W�>@�w7����'����;m'Nkzs��|�bF���.��)�h6��֟]H@��[9O�й#��}Z.�O�<+�/��p����`AR�㱐��:~����z�,�23|�w}<�&× �n�E"�L���MBJ G� E�a���j~��-CD�-�#�?�(�
:�i��>߅$�>��|ؐ�vY!�������7�����P�������k렽4kk�)U1�/}b�So��+������`H���`y=��k�ы�-6��IkLh����ht��$!������%��sј���]��u0̙�ص����Q�B����|�&iZ�`f�@�W���>�u���O�3Q3ƕz�k<����3�sj*w�O+D.�=H��R�����ے"�[K���Űg^�Ƨ%J�Wn���tyBW���헠��\-wu���]/Y��pdz����|YC��c��]@�:ﱆ;U����eMf��^"Y/rK欈_p��fށ��W5�n%q���Q�U-9p�k�D×+oQ)h�Tԋy^���Xq��a��w��wL�v�����ǳ�GR�"�H	q{	��}](Al�W����@44�٧"��u+Y�p{n�m:0�h�p��A�@����U�{ȫ���=f"�{���$l�:��=b��Sە�n�����פ�n��L�����=�ԹP�����m����Fۏ�Td���!U+��6��
K�W`!�1������a������ hu^�b֮6}_���Fwf�d��9��q��F�|���pi�ZѤupW�O�����e�9�6Ei��,�
Zi��R��)��ރ�j�b=�