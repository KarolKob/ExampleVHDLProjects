XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/rz��5v�	�>�����kPN����<h��p���8�M��f�"1��C��g8cM��q�C��G9��j��әZ�T-�v�Ⴁ�\$�Lu���J�Q]���J�WX�j.ʸ��qb�G�\z
���\k���?��6fX�׊���7,��^7��2�j|SJ3�T���)�F�#�^�޴�G#�E&�c�f`H��M6��P�g���c�/]rk�88�=N��lQ�O���Q����3��KǘlLfB�]�^ �7������\�W$<dB�Υ(��>�T?������t�S?�8�Ǘ��&��%��8`�ۥ.����YE��W���4]�vKD��A�S�'��%��/O��Mw��b�X��O��=bh]���W���a]g����G�����������_�;F��y�nH���6���_UY<��C�I��|��8�z��K-m�u
�|�ͽ�����J��~J����L�.vJ�=�2�ȑ<&�,�,��|��N �s��l���V����|��L�F�ص����s�*����V:PD6�d!�؜� Z�sB�z� ��_qЧ VP:e�s��Afr׷�DC������p�ˍ�'������ ����[�'��5Z����ۑ노(	�H��f����fir �&��4�;�h�����í�]7��^�Ӣ�p�V<Y(
�n�V=O�wxn`of� ��~�;�I�ѥp8��fg�7�o$~��s]���*�4�w#"��-%���XlxVHYEB    1bbd     580R�![�4o�S��A�O�P�L��B��SR��z1#݃M7�������g����>b
�v)
QW�y!r5��F���r�_1����1P��H�~dT1�v=�ڏUe �넓%u�d���An�?�sl��O���D%������(�4s���ӑ���O��<���T� ��WIB`P��AT5?�H����AI.v����Qҹ�� ��g�)7(t�봧�p��9�0j�-� p|��̹�yw�����V��G��#mr-�}�?=��~r܊&~y��y�2J����A|i'����sc�'����}���Gw|�Q	�O����D�LZ?[x���Ḍ�ќ��ˊ�+/}9Eۀm2�t���x�@�)��M��`�Q�N-Ss��׻v4��nPB�]����Gz�Hi���~RU���<д�4Җ���g#��u2����:�z�ݠ��Ke����]s](Q��,��g��o��$�y�+��������h��� :���k=�����s{�L�-����R�u�b��L�h�fG=*�#]$��m�x�OC�R��vO���d�L�(>��./�֘,~�v�l��~�P��lw[zo=��i0��}�kl�;	�����`��|���s�q���+-H<��ڰ���(w���d\[� �%�����S[�ȁiL[�S$n=5PT(�Y˷qs���|Bκ@x��A�W�f_[��3�.��`)J���7's��@W�#N!Q��@5z�H���Ѥ��ړ�=�69���H����1T)��Z�����O�ï{y^��/��c{1����kDl��!��$��V������,J���;�{�F�iF�Qz�(4����4�a @�2S.p�:ռ#�3�E��4q��̊��K���WM�	bj�Ռ����j��Kzزe�_|�7Y�7��]Y�r��cpx��Z�n���	kԋ�����%�<e�{W2��$�x�ZF�E�u@��B����
%xqd��Y&?��{�xbë���?�������Ֆҩ�>���&Y

�YY���h7�kU?�.�������e�зe]D��b�"`��C������f��U���mԭ"}4����Ҝ���!�� �sV Q�����u�=�o����{J���]vH_6b`:%��/SGW�5n~|8+��Jc�VV����d\�G7��*6��ǊI:%��L�]Zդ��a
�TheZ&#��q��l�e,�B�M�;9��Br��F�r�[X���X�
lYO���%�G��|�P�o��zO�,��dɾ�?�;������tF�6�Oy���9(���,���g���AP��K���d��ߋ���i�E��2)��hڒ`��K�����p��?� �z�c8��_��ƕ�t�-