XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ۉ�E�]��+%�R�B�����.b^:��ds^�G�����[���3�85i�X�ʟ�����G�|�i$?'`#��AMr����@��:x4�X�lY�/;��y��du3\�x��_�����D��/��&��d
]�11��4��o]��}~��뒅�4w���ZzE�\�J��ǉ7m
��ſ	�/#�����H^�fn�~�Png��;�"^��y������w]㕤��$������o�;tL���gQg	�I~����
����<;=����Gg7�@pZ���>�V���p!@iܿ-�+�j��(|At2�J���(}�l7ާ��/���	Y�Mu I����*��!�Y�@"�7h���g]U��}>P���>�̿���ʞt�Yc���
��?����y���]u�A]�z���0e�Mi���`����!��ͦѳ
^Fq�k$S9ઝ��vG �6'":�%���dK6�o�݃�G��`����v� EE���He��|��c��T��a��&���l�f����z_l�;{��h]�E�~Q�I����E<0f5��b+΁��ئ�2����9��a�N� ��FV���;����Gv��D�HsG\IAgB��mPn�QV����|�W#	�#�	0�<��>%Ǫ��8'�>%^_���(K�8ϒ�����k8�${�~���&uU�ca�٩�>��!�������h"�l�Q��ER���D ��9zz{=(��s���o=n����:��� 8XlxVHYEB    fa00    1a50#F �n_WMVk�l�i5�zz�|��7�o��M灇 ������2�(�~޽���*�Ww�ۚ�7y%�ʛL�L�S���p]�Lkh���@��Q��5�9ޠF̓�o̬`�W�P��]�cc�	�'�Rqw���oa�h�b�@g+R�Kl�H���̘P�d��>�/r�e�+�e�CsU��T�ĳ��&Id9�?҉�]�?���?Jb���_�P�UY�3�t`�����˘�������C��]�7�U�vOZ���0���ܿ#n�!p���x�����mm�K[y\7ms��t��z��M72&�3	���9���/M-� Z�r��;˶d����e�W��9����1ɷd�P��1N+����<�G_�
^]�� #:r������J#�g���� ߽$�9�w���ڦ�s!� ���ʑBN���j����6uv\w��Z T��ք�0�x]&��Q�vY6�p����D
m#>~B/�3��q�J#�_�a��-4dP0���U�,ˬG�m�]��罉F���1熌2�����F'"�'��d���*��c���G����y���,d���b5����Th�jv2{am�T=L��X3/
$��B�r �51�A���O�����>�V��:Gj��Dish)V�m����b�}s�k�5q[F:.�C��p��=̛d�@�� .���*��~ܪ�Oe�XƑ�݀�<�uҵ����˻��5�1l�u��P�5X�W�`-/O����BW��u}�Z��2��� L+�gЦث���z�vw��ۜ��9#C�2+�v��
���[=G]n��5 2]w����sx�Z��"�}~�1AO&��G?f�N�/�0�3 N<�N2�[�W�sl����i3��U��{'r��C��@��-�ހGP�d���>+�r��зNW�G��M#-KW��]�c9;ǭ_0Ǡ��#	����3�K���ESa�O{���N�o����C�rC�5�]��'R,Ss=t�%}*�Cr[(�4C��a�k3��� ���<2t3i�����߸�1[J}j����*��	�n��q-�t�`Pv��FQ��S�Ԣ=�G� �z{)7/l EE����.u�NyZR'Ŀ�L�b�*�q�����Q���.��5l��WÂ\.~�7�&#ϡG��j�+	A��t�6s�ȫu�������軦���"7�B��)i�*�ʢ�	 6L��O��ex��ZQ�.�c
,����`Y��v)�q�+�|^�J!�QP%��m'��V@��$�m��=�2��=�Z~�X����
�H�2���%����-_�S��vI��4}U!�S����,�£Aȝ���.��B*��R����&a��;@�����;��*��aK1-Ji��1�-��ܭp�0�a<��l�i@��.�@�#X�WBBC�F�Xn"0/_��rA`��c�u���]���,vʐ��W�6T�vV�3<_�Jo��>9b��[�����K>[�7�8\��v8�a�}Qs�Հ������ �zEI�ls��,�����p�8!\�D7m$��AsB��>���P��yV�@y5��_�ti��6f�'��+�����U"1t�8'5k����lho/�
\������}�t�8	��F�q���r������` Owdei��anc�Q��]���i�����ղ��6��DzA���o���0qB����Ӵ�U�E��?{:����סJ�9�gy�~��4xNi=a�Bp�*��]���p��ު�#��e>ȁ
U?!�#=I����ؖ&e��C<��o����Tj�Q�����Ԋ�WE:���@��z��J,�)E�ةV �4��D����mͶF�1�[5I�<��Q@:u^]��n�C�*�0��]'�.�m�6�T�~4����tU�.��Z�+��㯙�����1����0&�
�ɽ��}���j�"���~&s�hڀ���^
v iU«녅$��~��j8����Əxf��5��\�6W����ʪ�t�(-չ_+:�`٘?̎㲭Xd�W�n:�,j:�"��j�"N��
���xC�?d��]�zz�닆y0+�3v��i'�K��3\l��+����wv�4��*e]�{>�n��򧄨�����-)���=rU�2�6Tc��n�1!�x���mJ���N��%WT=�1�%��1R���L�ḣy�'>����A}cS8��@���|�潈؞���ᵓ����]�B�p.�Z�VA���GP$��EӞ|��f��af�m3F!]�Aɢ�j�W�,�P�n�Pʅ�H\����Q�k��h�&	�È�4�c��Hr�f�1�)%th-Õ@���&�Kj�>yn����-҅g�D+��;���Eh�5�Ԭ1%���[z����C>6Zw��tK{�l�x��C>��:T9J���Q�(�@��� w����N�Yu�-��� ��]��ֶ����W�c?ߦ9����������q�2��Z�{q0b�9����z���g��-��L$��e�j�@�<�b�I��1�|&qUa�l�W��=�͈'�Q(+bP�������tldx��@1��K-�մ@^FY^t�G���)m��]{����;���Il�X�v�(��#2�K��L0��Ʈ��P���z��u��KC>,J:�C��`C��ۑB�g�f�&��'�(KG��@& ?	����Rw��С	� .�w��򞀄:a����J�e�7��J?7��5��2�5C��U�u�i�75ј�b�*�+��5�0��.Ji�_�f8���:^ϓ A���L���0�zL��:W�3X�u/��AH�uQ@ץ�y��)n��?��g��2!��y&��C��g!]:���=ܶO5����K�m�`k�XL���<�[����ݏl#���[�6��!k��ћ����E���]��GSX��>������½���=b�Q���_o�~f8���C��K�u�˭QR����˄$����xR�45��*B��(`I*j���ksӦާ�P��������C���d��e�u������ts�v�!�W	��I �ݝ��z����biȒ�P�D�v�7D��_�\��>O��{ �-W&'�i��*����O��"?h��D'�W�N�2��|���K���v=��4ܥ����k�A8��g2)��!l����j�`!]�v�K�����R�.���E ��A�L��A�(ц����N��po:���	ݨqʺ񇴪R��`��>�����+�SZD&:�q3ֿ��3�� D�a�m
s�	�*�&�9��0�s��D�Y�T���k%�l,}CHD��2(6��9P��C
t�?&����������uG�<\��iBdeTO�(1�[�d8�uV�ӈ�L��Vl2�3�T������Ig�!��@.�d�oB8�g�Kg����d��Mw� ��GpsC@d;2;��A<�a���(��5���3��ѝݴ�A4p�$U7��9I�Z9�C����0un�bDwo�~����j~����'=-sA,StrrDH�B!��"�J@j�_Oc���C��4� � Z����ng�*�3��a�xڲ5����%e����Ł��Ț=;z ����.s��_�eCH��ڕ,P�?�~�a#�$��+U��x��"m�����l�	<��s}��Ԯ]/)}�GB��yFi�/'4q4���r�E��L�&�sl%�D��L�ZG	�z3ּ D�Ƃ�P�Aؔ��#q~��(kO��c�	'z1��/� 'ߜG˴|��BϽ�.K�V�m,�v�s��j�	
�k{Ќ���-����n��@j�*sK����0z5�y�9�;w�	��P���Ġ������xG�������0�lޗpV�� ���ť���z����U�aN�;{��wR�`n@�K���h=A��0��"�*�h�ػ�e����-��N�A�|�(����A���«X;���L&6�R����{�*�w܁� �T���B��,�V�a��Q���}�O�T]��䳝�����y�.���^s ������r�-L�>n�j �B,� _� O��% ���(�1�3X�J��;f�oc��V;@,BٿX�ZNr�Cy�;	B�m��j0;	�ɷ�2�4�L#EP�1�N麹I��Y��S]��=��ů�C�v׭�|�e֙E3�6&33�c6�ҌO	��Q�<3q{Vs7��yA�ESw���G�Hg����6��|SHr;�<Z�2���ª��G���쁜BZ��U�q*%�4i���w�K~�������ˤe��yۥ �B�+R7,@��أE���TXC�=o�Z&������zi����t\*5�0 �0�&"��7�5ʯ�{2��۶+�x��f��#FX�[���B&|@l���te�޾��4ssG��ʌ�RE�.��,��.P���|qYv x��rk�o�Y����Jm��D�91�@Eli��:�S���������o!6M2:Xk��9jS,
��<�r�4i\"���+���������B%�,���ϲ�d���g��{�L٣ă�kS�7o�K�!xԿ�C�cH�� Ưo�o|3-s���$�?�(�ŝ�$����Z�вLgH%
K�9��>��p�v%���SF��;~����E�@BV���a�"&Z��O���X�\���vI���Qz9�Y\�
/ x�1���������o���p�~;3pT� �b�� u�p/�*dFL���� ���t�h�x���@�"��OD,+�`cG�na�`ɗ_�#����ԈעH* �vA��f���i���znp�����X� B#U���3-���@�_� �i�u�\��}�"7­6�P���ʣk�``�Z�ѕ�Q���SU�v�2���0B)�t��d񛾆t��C$ H�/%�5>2��-ky�TN�lz-��7��������whܢ̓?���J}cp�e�b�$Wލ��}���F��V\S2��e���B�{�'8z
�e�8h�0E��c�@#�D��~��έ���lp�D�{/d5��B�b����Mû�C�������ȓ���� BF97[,�Z6�#8eۡ�%����b�����u �^�%:Ѽ�|�?x�V �4���0�g��;��A����2O���%�j�#�Ο+�U.�9cE4�QG8�m���~��_eC6��	1n�$�؜�kmx���h�8�K?a���/}�j�vR+��pRZ�{u���]�ӹ��\m�f�pa�����j���Šw��l
H'�/���بC�9���/����xD�D���D�DoWF�:!��W����8��[ӂf��CpA g�OQ��A���Q���ݓ�ތ�@���R+R���u3� ,O�[p�=��]�4��(7��B���Sc��ٸ��R�?�Z���9��SC�5B�OV�p�r	�yV�P䓺@��?�.L�$�^��+C#�*�ݻ��������Q6s��Ir��D��Aq�U������5	�}VR"w&c���כ���g��^Pթ��x�w����SĀ~CE��k�!n���ܮ+�m����!X�7���` +�+�I^�[�H��<�kE5�(Ly�؄�i��4���o2Z���g��NV2џB��D�>�j�68��"��dv���?��ʼ,zaUϋ��S"��n�тr��>�T>8��X���Ӂ�'��p޿Z(gv^�~K�� Fx*__�# V�0�l���&۵Sg���B�ڄ<YG�\��얚~�����Tpl���5�Dm�%M�[�,+��*�f9{"����Z?~g��#���hj��Ī���:��U>!��S�J�l�Km�y����A�0[���Mn��bwLa�#C�aRZPetb��j
���3����7f��P�5AI��H���Up��{.�_4�׾<�
��-Bтf�ʃg��a��̯����蠂i�{tH]%VEK��,�/�L^ɕ0��ۂu5�o�~A)<d6 v�N���޳g���R��ƨ:��+�:zW��F�
#�D�p�z�Ϥ�+`_k ��~y}(������?>34���=@I��dB��Z	F�>�����d\�5�e.b��;��!����ᩤ���~�s���`�#�mv|�&m�w	}�G�z����bi2�88�����-9=�k�l�Cg�Psl��%o�V�⮁S�������\󓕭sG��S���-��!X��5:� ݎ��"Oo�|C����<z�
�6��@�ٍ�^v�ڤ�^A/�jp:(B:pZpR�G�/S�c�^qo	�y�	��U���+D�*$��<�
i%*u�h�@f�՝9��e<��5�]�	��4^�S��@�Hu.��F�Z״+d E�^�Q�9V�Q��r8�&��r�u�����O�,ë��s>�418`ԕL��l�~�A#?E*�ވtaJn���$Q�H�,E�m�+B]a�1��4=��";�kOMR���}n�J������YU��͓3U!Y���!s���,r���-P�D�㫭87�)*�$*e�D~�[H��P0 ����8��j�=����g�h��jq��a�,O*���+�XlxVHYEB    a482     f40�7�^C��'[������L��?�D}�b
#��DIa'>K���V�3ؖP.{�E�F��FD���m��쯘HHF�Ki������ϋ�쐜y�j2�#��b�R���ܱ��U,�n5������e�8%�a��o'���E@�Vs��ePu��l?p`��_�R���'�&�i����	��Ė�$���?�Oύ7_I�w� K�ҋh��}s�Ǉ�J��-��ӂ,�s������$\�c�MJ%1(�r�:�7�L�薴y1W�Lkϔ�i��UG�Of������t5�2�� ��=�����"�o�_���ސq'��l.I{�K�/v@��g+b��Õ0q�.*щ��q%�AX�͇s�=�tG'�&@��'�{�� dS13�-�����X/!�c�(�$��n�X�T<M�s�Ϗ���U���i$+�-}�PH�:sKInΚ�*`1@�G}�z/J�e�;���|���6.���� ���re^G�4�+����yU�Q�C���f�D>�di���]��ƹ1g�qΪ��̦YS{ޞw�vI����;R[_���%� ?$�H��5յi����$0���\�7e*4��!��
1�P<�-ERW�}�A9����0E��׾b���z���F8��*r�^q�ʇ�4�'gk����D�ަ�0*����r�G��ш�-O7.o4N�'P����!~�xC".Dq_k	�Æ^V�*+�U��';wox���KY�θ#��v0�)M��w�H�g��z�j'!ce}�E�[�b}�$t�]1�<-��1��v����,�]T2m�i�$+?�N�� ���.I�O�!���3�JS��NPa%>?y�˹�Jսe˝c��`�A�!o*���+��Ю_ #7���$���}@��k<F��K�	�"^O;�#43ƺ���i#�MЬUreKy\|h�A�������]o�-����\�v���&8���1�pA�j��	�B;t'iH��ChQ3%Չ��g�X�����Ǚ���V�i䂵�'l`Z �ּ��0�
��ⴱ�]|���h��o�R\l�e��c�<�R=�����$r5$)������������έ�����=�O[>U<�&�ɍ`{,7'2(Ð������@�f�m��ҭ9�H�\����Ecٛ�˂�<�s�eaz!����q�b��~��G���{w�T&�:i�(��3�Z[����:�Gw�(q��jm���x�h��%n�B4�Gw$����[����K9��o����,�!aֻ��g�+��%��ݥ���I�h�v��o6&�[��)��� cf��{�Iy.c��[��$�m���j?�zh>�1�ȶ��1ي����"�i����u�0>JP�%�B��w�
?2cZ2B�%�^c���~��)��(i�O�qE����pn���s٘N�:��6�f���V��1��Q�w���2�dT�:U�7�,�ݘ$����4H<��p~~w5R�(Zk�SE��k��94���rT�f�DdK�3+���5�+��y�p�2&��?9�&��z�l�Mw��(�
G��*t0����p(�L}��k���Q͊��n�O��|ؙ�?��ߎ$FV��!V������0E ��_�`&�jP	G��;R���@�-�(���n`�S�X���J�%C���2���<����y�/g�w�ik�$D$�yg�eT�N�wb���2�eU�� �g2�uh�"����[mgh�3�H���+^�p�/��������;15.�v�;�N���j����o�bj���Ac~��-�}����DAV̶�-Rԏ�AϜ�ӄ�!�z,(N�A1 ̷�����i�Z��Xt@S��N�w��В��g��)B��ގ	��W�)�-��J�h Qx��?r���6��v�N������fFū�ʕL2��}�ӈ�
u#�`�DɇW?;/vE	`�E��޼�s�˕�xg ��=�r7+!�n�$�a��`�f����9B}YM���'��K�����[K)?��a"��.D@�< V��4�d2���z�<>��x�ѯ������¤�j���!m�q��"�s=t�ݗ���Lw�����u�����+1"N���'�s��^7�l/tΔ�e��r�ҋ[ �qT#�N ?I��q��䭝�vkH�MI�ktE/_�M��'��u����d�z�F�.Y4�U3d$����J�,�;��������-ӿ\�l���\�1�Q��+=ާT��4qڬɂ��,�҃d퉋~��9��=(!lr�)��7m�J�)��c�!�m/��,~J�ֻ��V���w��C��˷����SĜ2@�w��
=�&�!b���^^�s��]���W�QZ���k�m�$@܏��^
�H����@�*��B�|EFh��I���Ԟ���P��B��k��]Cʲ�x���6�}�o���Յ{o�/�6lÝ�쪻���coP?�'�Eí�i6����4G�|�!JL�W7��4G��hTޏi~U3���.z���gj(�xS�Yk��":l�BD|Am�;"Z�Tz�Zg 4iz@�$���|�E����24�=���2����� ���
��{}��Ա�\�JV��z���ۇ`x�[�e�/���ca��>�p�:�h�;Q�X���X4#P!��f'�/��9�˓�*����f߁?��N�-m.�;)*�<o;�p����ѕ�E��'�5��[�,){��K[�͹M�yx���Ӌ�y3������wc��r�.�ۇ�[L��@���]|�"�/��$gj�^�����4D���~8����f�BˊN�H����x��㚄���~5њ�O�����)*��B��y� ���z!�����n������J�)�{��A>�m�N�v0X�%Ɖ�l�S���sr�/$[�q����iN_h��g�?��+x�,j�� �:�*��pj�k��������X�I�cǶ����wn]��~r\}^�O_��b�8$�QV�fE�.|�9&������=x�Qo�nO��&5"��6�G�Npn�'�G�^ �~��^�HV��րț�rg;�|�,��)�]��c�A�%1;,�Cq�z>�����1�ٯ@�r�Q�i�� �9Fe]�1|�Tvt�8�L�����(���ׁ�#@^@@$�wMGo�-ҪQ3Jda�ou@m;nk�Н��6w��3S���XЬT]��G��w��W���V|a�;�^#^�c�bB&��!1��Ėŋ���]�,
2TEÚ�49TiCEu	xz�E�pϨEo���n�Ff���;N�LJK��VZ�[�i
ڮp(�َ������n�>z�[�ΞN��d{>���ƫpf�cA�]X�}z��4T��w�%�z�A����0<[���/b(�e?4M��J��q4���گ�C���ǂ�s�V�%�A=�H����W��]���b�X��p޵9�D�Z(��r��<	cM�MgD�|���\��B�RQ�����t�uAց�A�V��=�*�B4�U��B�(X�b���9���=�5�ge��-�_c ���q�վ�}z���25���=]��}S �`����vM��X��G�(1��c���v���z���Y�	�mo4d8۵��?�e�)��`1[�F5���2��-�̎j�yVc�U�N����l����\M�4z���)x�(�3�z�?�$C����X��Db��QQ;���H�L��-5�������4�dT%���>a�Z#Ǐܡa7�%��J%�Z}���XjU�+�a�(������.Jj��e{�Y�^��龟���O�97>#RW��A6*/��