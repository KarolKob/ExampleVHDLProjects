XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y��Ë�Й�� 2�h��k���C��m!ܘV����M�J.�W�x��gA��ޕ���Oe�Q`vc���������黬�֞N�����2��W�)����0��ӻ�r���G����L�����,R?2$�[��Q6�/�{vH�����z��C�X0w���x��{�e����Wc�����MKSΥ<|�#���\�?�����#s+q��l&�ž�'766MM�\�zY�2��V�`�5Y/|51y�l3���o�<�,�j2��W`�R��Tʘ5�_��so<L��,[7���F(���y-�Q�q��a�d�h�1��6�",W�Be�韉�_@_�K�FS���W�2��=��5Ǟ�G�(�Y��f���L���g��)|(❦��i��߯b�D���1z�(�
k��zJ)ڀK��YUO@0Q���\l�cf��v���`Y���a4����҆��x����S�Ա�J�u�mˉ]]댥§�J3��،���hI�^��3>�7��?���6a�p���ę����u�Ⱥ�qX�P__>d�v]��E�iYE�
�����7E{{+6�)��[||4̠��U��Yή��oL�Cvm�=��d�_�Kr�>DT�/�y5�W��:��Âڲf��s%%ې�ǉ=xTpZw0|�t�ǥ��ȰT9؊���C˷�����9*G���]�ܝVJ����P$ҵ$fXX��u��������D.LՏ��͟ ���S%1w՗,�eY��Q�XlxVHYEB    2864     9c0�icC�Dq�ʻ��4��$���8٭�\㌪iS��0B���3�y[�c�ܻ��bFk3ѐ����~1(��1�*ʈ���(�lۀ������� ���-����ӎp]��������V�-E���ԃ��2�w�t������\z{/����>���[Օ^#�Bn*��{Ɏ���k�[�S���0�Y������Vt�s�?Ll/�@~�N�;���E��T�؆�ې�Du�,6j��xg iQ]8@��y�a;�"�VpM	ߋ�,�_�u��Dc �ӣ�x�uۚ��/`��S��B�f�z�>���M2��I�#XZ�k2��O��?x`Ն�p&Ѻ=���@MI��˫p#W����P�̉U��T��rr�8hk�եuz�B��Mc��h}��P��(_ߐ�Pgp ��P����乊,"[����َ�1�b ����}��vk�-�)2�6Z�oCp����kUۑ�
�ro ��oP�B�b-w�;��fL(�Q3��"��Y���Q/s����d��:]�F<�"Ty�{.k�Hu���q���z믧��wV���"
D.~䁚�$<^�Ǻ�|�d�d��Ж�	�6���G\�eF�:��+���U�uI�*NAЙ���8��1(�'�H�9�̯�&c�2;�5�(����ܕphx�$����D��l;.�I.n��U�-�Eˀ���R^������D���塲u!��2U���Ӻ@f������U�y�	�����U�#��W8����)�XT{���Q<'�����#�"|Xr.�k�V��-��zO�(����Z����h*k��km[�4FPU��	`ʹF,�w@�W��]���46��sKfb���
l`�KR_p�.��^���5^5��x"�>� M�Z�g<y�5d��M�Ѭc��6�/
��L����^?���y�)o�!�*�m���pDʅQv3AnϚ݉�}M���y*
@��SfDs��~eA_4˱�l{/��|���|�U����dU(���5�լ�V��k�	�W��?C�f�dy~0����d�j��,�L >AR���Z�s� -HHo=�w�3R�;y��D�`�T0)R�`��ym|���~���"m�����*�V�)jmuz��#�>¹��L��{|c���X�D�m�Su�M��Gj`" ُ[z~��hy�7y^}��A-a��v��b�-�mЀ'����S�.@Q&�C�=d�FNuЌM�iaN����ݜ�rPBL����U�!5�M���P��#�!��w&�7b��ȿuT�S�)�G1(x�����knj��JP\@j�ݝ%^P��ר����J*�D�hM���ܨ#`����$��]'W�t �B�d����-���rxa�v������'3�#���s�`��Ĺ;�X�Y}TC��s:�������,CP�:n�E��q�<�����������	>o,狈?��0[n`��*�D\y'n�����p�6���G��n�>�!j�!�9&><|��	�p�1|�%1'�9�Laޭ�Y�<9x�M̓I;���=��?�%�-b�y�uC�Ρ./R�t'���'!t��k�<����(iU@��-�wfR�	�����_|�X���<y��V/g� h�[��7:m��ؼ�j���pJ .�j�����m���0b�|�U���<?��IC,�8hl ��-'{Έ*��$�n���Ϧ����8��r!>Hm����ޏ�g�E��Yn�O�jͬļy�.�џj��M�D/}�߾�����ٸ�K�Vh���.7����gUP�E�Wu�m���Y�܅��J"�����:���J��8^�B+�	�-EA�wv��S�;�Wc����W��s^2�ւ�㌹]F�0.�^|*�*�7�߹q�kҷ��&l��m��Ҟ���Ǽ\����w��z�-��&�6E��t~����n4�º;P��?�+B��K&0XE2�H3�+�0�g�E�x-y��w����x��Ƨ����p�>�o�?�?��)J6���R��k�>��P�0����s7��fTV��E�"�r��)�پDtE��f_WtmޟHwK���g���7H+��t�I.ǨZ{G�kX\!�:Q���V��gW@�Sn\Փ���ř�S�_�J��E�K(ʫl�e�-,��/��9����
�b-&�	��|�W1�C�E��:]�b9���p��~,�D^l{���Ru'�����z���٨���u����}$7���",^�iTZf�����;��Lš^B���'�]4��M�����Q`�x9�:�%����[;��k�cNؼ�ʹ���L,�l�,�I���ADu����|����� ��TR�~�%	l;�"VȽ����d�o2�Z{��	��4��(�){��!��l����B������ո^U����s�-% o^�c�U��fe��V�Mm�fn��:�'