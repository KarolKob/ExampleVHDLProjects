XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���H�ΤB�[��)����l�G�Āj-I?��̵��yj"�-nB�Y�̀�;1C-sܝR4V��A���Ū]3�K�ĉrCm�+��0;��n�Yj;�μ�\��-�E�].��:�q�ՠ�T����$�,���f���Wf>����#��|��쮊�M@��sͮ0E�X�̄ǩ$����O�ۈ���[LV3Y�c�K�3��p.������#50�U�&lI�;��	�>��-�� ��څ��cl��]��
/=&��b>��{~%�/	]�N"lB�,H�ۍ�B���
��7���f�O��u���u��Qv���&<�v�fݑ-;;�*�b�A�����(r�X9�N�L
ɿj�'�q������=�INFVv ���3��h7A>��N8��Gyܢ�@�A�7�+��dK��
��7KB����fMvQ�,�kw3U�V��c{��]�%�{5�+���KU�!t
�EHj$:�M�E�5��pH���I)m��?Ș_���.��4�J:�w6}�'W�;�R�P<.��}�}e���}e�E��R�{#uq��tHd�q^[nxι��:��5�iIk�[����$o���vl#t8ތ��j��3���A���`��)mD��r������5SrYY5�k�Q;�i�Z��p�Ti�<���w�Q�{��<����D���������&�f��;�X�X';7t�!���ͱ�B��ޔmVF�m���tO��d���Ք	���]�Aap�t
�����'ՋG;��XlxVHYEB     ab5     420�gC�\w�N-���}��g�/-�Y���#��q�xJq�E��8�ذh3�;��;,�j8dm�������x)^�8pj�^��3�LM��D&D�$��J��Ҋp�/ݛX�*�s��QE6�i`ழ���bp�H@f�{�~o~z�LwL�[ה8�%	�#�?\�/i��:e���)mS��ʣy���<r����nUDk�?:c؄����Ֆ�����7�ލ����|9�����!$�H�6B��}�$��JI}^���֧��j	lK���L|�H(�tښ��4�SE���ne?o�P�_���P�Ltp����ј�|���K�7�;"�h��.����
Tp%|z1��t���tG�4�e8�=Up����z2�x//j������Z�u��HJv/R�����\��&����Nձ"��;V�Qg�mu(ԥm��~N�����4��ӕ��R7Y����Ư�=�?�F��cҢ�A���f��r�����d��F�eW����{�*|����n	��VB�rZ���F�j��KV�*e�v�/U�������;�T�z�e�R��=�A	����ϒ��@�l�?�+�P��5�{��Kf%�%��Dox d۷)���E:.�mem�ZG5!첛�%�9><��"�y�F㱀�$k�x8������ݚԶ�|��M�G2�i�_��G]�EL�OF߉��э���;�U���WDPw��89� �u>#@,�(�&u'�x3-Mr��8q��G�@p$�v>Ϡ/�Lg��Y����1�N���������ƪA�(E1)C�o��?<7��=1 b��"� �����/�	�خ�=��S������6�6�߲�4����tt*�6�ab��iM::�`��	����Y�N���\�4[.����m=cQ���&9�������~��/����E,��f��xx�h1o1l�X��e΍��g�?��7�er�l��]r"[�MBF?�8�
���nH��=�R���G�WW$�C�4X庽���q ��D��my�kʌ���X�