XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� hZQ��54S:-�1�n$�T�֖@b�;"�օ�W�� �
�S�W��[,��[Dݓ�v�(t�����2bz��G{6.��*��Nd��HG��=wb��K����i��2u3����y�x8�ޢ��m�/O8~�]�KV���,f��F
���~I��n'z�~ d��a��S�3�e���~w�Ϫ�weNv�^3(�~��~��q/'��,b��#���c�+V���K�4|�&]��Y�X�[#�fƆ�}�`PkqK�A���x�4�	��>_α�_v�۱2Jd2�E��0ۨ�.YK��������R*�*˕�=���]��P���%B��b�X8�H4f;%��CPӤ����8���r��������knM��m�	�g�v��G3��(��9��u�uֶ�y�{���3�5Q.����"-&��W�Uq�"i�A2�^\�zQ�n.��H�
>��ޅ�;O��B�3� g�솔�������>�(A�4k}���Vr�eG4�8��ܡ`V��&�!,C�j� ���Ǉ�_����z���s������[���O
9�)���pGȏSEm�t�a�Ĝ�H�M���Im* QH��ڝ]YI6�MN���!$AV:��
f�z��DO��5(�_^�Ⳓ%0�E� �E��$�Z����p7�Z ����[�j�n����}ݜu�Z3f�.�΍�js�ߥ�.�l���6�S��V�TW��Ӎ��E�CE�`kdε#��G2ڦ�ӻ�u����k�O@�J�!X�XlxVHYEB     b05     370l��JB��S��� ��ۜO�@�T�%��|�nh<�`�{�C;p�E�~?�T>�1��lBh[�t�X�:T�c����
�� �Z�:S��nSa�]�~��Z������
xx
�O�M%H�t�
6__n$�ILN��Ƅ�U��3���@G�Y�	%���1���Væ����=s$�"swado��ҾQm�� �3z}�
�oF��q��O��<�6�zF&�5μ��
]��w&V*���Q���U=_��T{4{�����n�c���w7@��S�e{�L����� ��l4�5ˋ�E�6D')0�6��G@�h��x�}Y�J9�n�Rƛw=�o�.��r��W8b�vJ�Bw,ia��\_�Zp�&B�|"=�aB���C/�OFD���;�/|����`�z�"#��'�,�|6$�FŲ�䉑��K�כ�<k㴑�W������G�p�|)��|�7 2���)F��"�r��6Z9��m4���g��rz>�U���t��!wb�9D"�P9�7| yK��Ggd���:������*����vv��߄f�l�X��j��o[e^K�NzoO�͑𳈘m8��.��'W�s�w/�{W@�w�`���N��Z�v	��� v~�ҲL�%���b�R��+Z�� ꒃ{#T�$g,Lj$�R�H�Ԭ¡�6���h�hO�>b�s#���ޝT_�;
�Mc j���6�()c���'�i>gE�<ɱ���FG,��p���.�AOܥ�W�����/��1�ҥ�S>fv���_ l�\rgǇ�"���yV�gM��ӹ�Um����?�ְؚ�fs���;c�뗋�Y�m.�Wʿgf&�P�dw#��Y