XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oE��:\}�w鎟.���E�v�±
\���'���t�꺥�m:Wk��.@
اC4��ǲH���;(�۳>( ���T������e���
��'T��o�f!0ڸ8:�'I4x�V�|�7�G��(�ݨ���KQ1L�acf�L�X�{o����xDl��ì��j�5ǻ�h���'e�0o��;�r_�Z-�}p��ް��Yx����j�K�~ov�[�iO���m�� �+^�נ��aN?��>z���Z0k�8ԋ�p�ǥ40��}S9�?)���Q��=,E������L2����2�����a�?�6d��6��)� 6`Z� ѷJTcn8�����Jl�ɒ��5����J�9�+��vB$aw`O�5���{��U�3��;����JG�oX_=̋���B�W�2Jf�����D)(�"$I^��k�s����S���a��ۤKx�z�J�^Nx�͒o3���C�1Y7'p�^�$��3� �������3�7ܸn�ʥ&��֌�i�دmkq�X#��eL4n�eM������䡅���CT���o���-����)��v��#�yz檥q�p,+��@��^��W���"<q����ɛW\}��$�>x��-��H��G�����C���AZZ��L��5���Db�'B�^;��?��U��B��lX�FG�EQi)��֒���(ˎI?mM\ʅM��Grv��)1��\�P���݅�� �uб�U�W��3<��XlxVHYEB     7b8     2a0_z�F~?�v�F��#5����GX��PQg'���]yS}��c�ib!�$A6�J�H��z�}�~�{I͹�55��T��*�m��A.�CwIX�y{�lBN����O��H�C���3~���.�;��ƿK�ŨgbѢv�jj�M����!��������|�
��IQ�����w�ճ�)$�P�7����H�QRO%��)t",�1v8�,��d�=�_S�q��F�4����7���֎a�Ԥc/ ��<�d>Л�� ,�E�m� ,az�D֮�WbQ*��2��wv����{SY����9(��Q��\"R7���Rz��]���TWvUn��ԧo��+n1Ė������I��lI��8�	d��߻X|�wd+��e�����+3�w�5�`$�E�	10GMկ��l��#��/�1���vӜi�[�UP��Y#wd��z��r�p����QR�c:�һ44k�"yet�y�fV�wi��6ݾv��G]���5zzQ&�JrV�>Xj��o��)��C��KP���h�杵|ߩ%�7}�? �֟���p��|��%D<	l�Iw�^���X9%�A�m�:ި̫��p�����1�St��n��0�{�	R5�9��T�-[䘓�Ӓ[dZ-^~@�x�چ��;�㰕K�G���_M�;�n�L�