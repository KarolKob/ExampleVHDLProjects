XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���QUM�J3,n.m+����d��� ov�@뭁8�rò�$���Gve�������	ch�~�2v̮b:��7�F�[;���ӹ2��o��F��t��c��pV@}�9�6�D텘�R^O��^��O��\RA�#(�ͨ�5�7��B^��ӹ	L��͐)��pն
���貿[��^��%#�T�%a�$����FI~7=j� nyW�,���Z3���P��#=`��JM-@^�NO��q�ɪ܌�|��;���sm&���-�wC�������٣�[����x0��$�9�2��a�stG� \P�ɏ��u��x�Tw�4�ڋ��k��M�}�_M��77�V�2�'�Nw�׵��HP�V�4���D��\�����N��O�,�v.��LB��h�o�����v�����AƢ|�5�Ӳ U?z0
,��*��L�DIU,����"�&��
�b;�ްCf�a_,U@��<��	��jm���荝5X�bW�Q¨R^���͸���9SKe�U̙��Z��B���ݠ�/��V�*���W��|�l�q�����S�Hm���涾���3�������e_%��2�k��x�����U���F��A\��Ȣ�_R}O<��0�6�f�^��p/�L�D��fĥM�N�%�w3 }�<�z|c��v"
��� .��/bM� ����txE 1V��>�h�`�MQ`��uJ��[��)l��D�
�]Gqg%3J�(gg�p���N������XlxVHYEB    2d5f     800�t��2Y�1+�ݡ���3v�����-X\i"쪏J���qǙ���6�� �����|Hb$�)@(���Q�"wG��ƅ�Td�P� G@Q�k��C��p1�I^���c�B��I���g4h����Zf9�ó{M|w�uO8������K�L��Y��I�p�FD�Y.���щE0���e�wz�V��[�^Ix�T�:�xߧ5�Fn����
ke�b1�k=y��w���T�-=�d�K��2�G'Վ��%�3JDD��S:tM?��M��T)�#��晡�ܖ��dh�,��e��?Nb���q�ANN�gF书�At�U�
��o|�5���_��,����H�C��x|�������8�R�E� Z�bɨ6L���2N�.Eo�V�ÎP��0q����~�"���M����T;��R�X�j]�a�n�yP1����%�rH�D�u��\���B[(�F�?s�P=|(S}�ƈ%5w��1dPoB���_f~�G�~O�Mp|��6'LC���{~�y��:� 1!499�q�\�4HG=�i����E:��L"Kq���*m�k���l��KO]d5O���>*��i2��d�V���f4�JNe��
0!� ���|�їy5L.��o'�k��;�r�D��EM��H�?�7���"���@Z������~c���H������7T��nJm�`v��ߍ=��~x�!M� w�A L��P7	���K�#� ��lb���?ae�}:��)b��~�O��| �y�
��mc�J�D+�$��7'l�ִBi��e�K��`і`�э
�R�g�D� fw�� ��*���:�6�e�rE|Kƒ��=I�'dY�bC�Nf�r���o`r��;(=�6��Cş�O��Ƴ(;>���V�,-ko`o]��o�� xz�ޱ0�ja��A�y%�%8�wՌz�)ʇhz�X���4�N񶟏�{.�)qҗ%0�*��$8�.�g#�2���oT��?gHY
_ڼ��S4Bߦ��Ǉ���5�<�٣�=��-��Ү��%��kI���^-S�+D�=�����Y�|���]��?�cnx��nl��a�2Q5��[d)`��&���DV��3�;E�s.���+ݡv������Ή�g`��~0��[q��N��;��0�琑���Ί�E�(Q���j���䱙Ta���}g��:�0�h?��n��.�h�DLzE0^������� �u�U�-��i$eɱP�W Ur����j�5(R�R�w�G����7`3%]%6A��
���h���ס��T#dd��h��E�D���1�C��MZ����2˟*�T� �	�+z�ڳQ��3�fa�����K����\������wѶ�r�Q�ZQ��	�G��Y޻�N�;G�����G.Ƀ.�5��1�m��e�BW�׉��,ZE���zo�yÃ%g��e��a�]M�!1�!%Q�.M�����N�K(D�����m�&*�S]Ats�EI��I��Y3�,o��1�I?$@۟�Aql{��lTU���ϼD���Yp�����",N���]�gKV)6��A��Tօ���q9�w��Z��w�T�����$O�BK�yޚdg�ΛT���B{�=c\�In�M�@�˷c���ժ�1d�)n��R#k�`��(�l=�`J৻xbx����x�b����r�����h��x���:�Ю��g���p��:�w�m�3�`�����Z��OW�gZk;{��z�!���nC���Ei�1Y[���3S=����)X�q%�38F'I�%�y럐I������f�/��,�������@�Z������j[|��*c$r��9�Аf�lDP��?�����f��L��C� �$���?�~FSS�"w��.^��V���Ӫ���fx&�ecR7���X�S�[ԣo� vg�۲�qy�
���Zޅ����N��� ^r��"������͚Nw�gp{�|S�~�"*N�_�x�ղ�^�D,�wY% �@��'���H�T��ĉ�y����`-yp{ˢ