XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X1�T���u���v�}a��ڠ�i_�CL������� �`]�ůq�;J�+݋��!��?΁E�Xu'I�sl�~q�F� �Ǭ�*Qj�mBh�q���D����?�3�5��������kګ��Q�Y`lN�x�L�=�=܊��{g�Ãsn��:�c�f������5�5�PK��Dq�`�����[�+\�8��}n},l���[8c�ˢ��/�\u��:�y�7Cr �Eh;S?Lp%|��8�Z�$d�'����0x(��;�6ɰ����Lk�XN���t���F��chv+��о����^�7�^��M���j�ư��jF���+�V�_���,�{�?����t���3ؙ7��V�X��օG��`�hj��|c6l�ܳ���ի��l鞫���e���B�fQ���'�{����^������y�OK���2�^���ޒ������ZxAE��#��V������R��[��1�;�'*}��QG
w��.��������u"ߓUgٗ��?���]>�� f�q��$�lՖ�K�9D��W�"�h�O��ظ���sA�����S��x1>�}^���k(�g彫��Ė�bC�N:��i���S�f@������cf�c���9Jp�k���C���r)Řk�3ro�SL��h�w�Z�&��y}�ͫ���)Lv	�|��iMg����-�B��Rf��mjf��P�������l*s ��xB�0��Eثd����� t??XlxVHYEB    cc3b    16b0FZ��h�w�ϒ��
�.��?�ʪ\m�_��(�+f�h�J�њ���#��]v�7)��ל�Ꮄ�^+���� ~�XeH�C)��js����&M��-Vn�~���$o�*1��$�f�����Zi�cFg{�H�������з���J�
��?��Y�{�rQ�I�'�M�*����M�j�s��>cá���$�vda O�k�
�d���m�Ƒ5�
�z�FFK���Q�zI�������(M��1E��K���[ã{q 88;}������[��@��' T�y_�/�8����N=�s�8M�*�v\X�8b���)R�
{ �PHZ��=svĎ��� �k��V�"�T.�B� ��B_�k68�"&4f�k5D ;!���C�鰟¦�u��y�б��$���Eq�O8Qh��$Yd�FQr�y�Q�;
S�ޱ����=�(+Nɸ���@[�<*�M��6��&B�L�vx�Q�c�Сx�.���Gv�H'��m�UOg�N�>VPm�T��k�R�8HQ���	IozP���㠮����b��zr"�+��Cu���1�J�ˣK�nP3h����OxK�mr�!�o����*�,���I��٘����/��$(��8$S𩖉հŽ�gTWǨO�<��-�A���ihF=@p��&m��?<@l��m�Qb�d����|�S�OY�3 #���'��m�>� ���PL>Mы lL���C�����A�� �Xqf��0�7��bL�@S�DPsc?�<�����6�����<�a��ֶ@���?�&���tCT躒���x�pN�k�����v8RŰ�,�����0}?q�M5�G������$�[��]��F�D*�J*�(;#S+Bnlҥ�o#���
�^;�g+t7>��>�nVg�*���}�?I��\�D=<�	��#X������v�{/�S
��(A1�	�Hۼ����zU�]S�/ ek�}��G��4Y��\�3|�Z� ��)�%����I)5��ړ�MJ5���*>Q���\������%���;��:���NՂ�UAM̔z�&��(\?��IZ�҇*�Ď��<�f(�����Ԛ�.qP�x�O�z.%��2��d訉�3}ǃNa�?��'��6z��ci���e�:;�p%�H�H� 'Z���Gb���+���T֦�ڊ6��)qF�vܱ��ɰI��w����5�"�1&��QH<͠�Bk��+1��ۏW��#�����z�H�l��l��}��>W�U�M�Ҩ5��'����֨��5g&�Zl��m��V�٧/��)%M�m`I��6%�e�V�=����<��O��;��+�/Yr�w�̝���x%��N:����H4���:V�k��@}�! F2�N�+�Jn��|�˟v�=�l�J���H7B�k#Y��q��u����f�y�\�5��EP��?Nk��˫[�g׵
h��n�c
ٿ����I��V~�1ƿ�����X�G�R���tB��&ir�W����Զ�8�z9�P�t<4����V�=�#0z]�-�����UK�V�>%~�P�;��
z���+�0�^xb.jq�e��靍��ȇ?�γb��(��l�@1	_Jg��8���i�ϧ&)��Җ=��A�&��V�=�^��l��֝�S)�ahK�������s2��@J���l�n;��Z*g�D���8b�q���A*v/P�'���U���h8���/���pL�緲�Ϧ0w�vI!#�r�k���N^�[�sn�� r�D��k!����ܭ�<�����ţ=1��/�mA3�RAӧ� #�M�'���[�����e{�raD<�^.��ۀ1U�,�ݰL��/>�F�O=�����z,Gy��$̷�.���n�͸P	m���z���~"�ȥ�oG�c &�x�H�DD&�}���0�\�S��99�N��|?��=!V$�t�>�4�F�������{�b����o��Y}�ҥ	�/H�p��I?�$|�aC�>�Dpk���$.YP.��u5D�k�&%_0��2B��,��CPZ�P+����&��8�3�Y�"E����|�~ح�do������$�WlK�����	q8���9�<V�mtI��%o�3�� ����
��/y�"E��J��Ѿ�)�����)5ߨ4���L����c�-,��P�#v���>:5�d��
'|Q� NW���[�=��RYU�م�E�o+L���9�O�����0�J�����)���6G9�,w���mt�J�#��7�n�],I�u"DƿZ���]�\�V�6�hz�o:W��@⻬��P~Չ�#�?  �֛�<�pڻ��PN�Gݯ.�*�=�$�Z~%��j�`�������,\6�����*7���/��W_&���st�5�rd��C�$*1S+k\Ai�9f֏�c�l���u÷�¢�C~��VI����l>PHȎ���Б�Dk��L��T�f�W���)e�"Ƴ�c��<_GW/�>Q5�-��?�C�b�6��	��?_vs���c���SzP �֖��
4��(ʯ���*Y	g̪i��>�����p�R�Ґ˞l���?l���LԦ�"j�`�TNo�Vv�b���2ᐁ�2����5[��l�d�v�^V�K@I�DAT��%��>e�+�E+�ڵ�jZ *�eK����/��6p_���u���7Vח,�,'ߴ����r]���2~�� &������7p�_�M5R��F�^TXsa�]n.�~���?D%
;W7/�'s�k���Zm��@1?�b��c���z83�+mJp��C �Ys�wu D�%T�`lnVK�������'�?�)/Y�.�j_��ʶ����g��;�>��⣼ڕ��e`/#!MU"Z�LUn��T`��R���ܽ�FP���k�b.�햿��3a+uU	C ��1��V�!��)�	I��h�?�݉A�h����VPV	�GU��I#I�Ȓ
�I�Jg�.��$����VQgf@n,�`8]!zvB�8!�y�"�ٚ�c�>���i���H@ fO��Ji�;���4ͮ�c������J�E��:�ۂ��潇���A�Q�~�L�ٹ;+�aI��2��$�B8�gs����$���ٖ��,h�cj9�=��цk�,#�|+g�vn����椷7�bx�9??w�Q}/x�k��9M��YÞ�U����%�*��1;�5{w4��6����#18�j����X��`�۔*5*���<p"��֕EOWX�_�_���a��_����qc�fJe�t���Ec.���Ɖ8����v�Նc{�	��ː
��9K.��{C�Qp�a7�����S�]�ea �ip'P��|<W�$y�&�ơ �(Qv���0H�I�g�m��NG���� ��C�T8\퟇�����pm=
�	vk�2�z{�J�Y���ԉ�G�#�h�w �
AI7k/'A��qMV��'���U��|sʞ���w�󭙷D�u�FtgF����^�a��(E"��s��ʓ{�:�H�Kv�i\��w��	���l�,`o��vYޓ�v�O>����L/p:�$�@�}�&��B�5C�E.Uf�9�M6�#�����i=c�K���!������!U�y{���CK���y�ֳ��N_Un�vI��/��UV��"�.s;w�Ac���c��#1���~-�9ȿ�t���#o��*:��[�鳉�X��P��&�o�� SNg<&��P�{��B>��;�
�Jc�,�Κ������Tm$���.w��������9~
	_`cr������iZ�M�9e����������H���\�>��}V����K��+�����VzL~�W�X�)׿��z����M�@F���{��-�,7C��uf�f��{�C6(΁������G� �NL!@�z�C�F��L�X}�[�tLv��E�JE�f%n�h�Rw�k �c�
}�C�e�[�{��b��hO�-�x��$��Ke2F`s��I���#ă�:^97�!ճd��׵�`�,�藹�Es	9����l�?���s�n��C(_
ʬ^D3����J��[6ſ��F��7]���]�X-��9���YD���`s&v�6�:��Q�LW�L�X.���ܜ	�Y+l��|8"�-���1�>�$���wvU7�k6�P]���<o ��E~�K\1�{B�:��$�Wc)8.;*�Э���s�{ P����-0-�Nu����o�����O���5x��_�+�E�����F��b[��ҭ�~j���~]��I)y�v�p��{xW��PWGGF�C�I��]�s�3F����S}#Yʖ?6@�X-��O=$�7���������-�=|_�\�T�6� ��)ac�P�|���w���?-�k�7�D*�U���~�|���5h�w�2%4�+�����_�S���sXu(t�"
�?��byx;���{�en��=0��e�:�$Pp���0"�NO������Mm��e�c�:�گ'͖\�4DY��Y�>�W���ԩPѪ�2�c��J<��71���`k�iJ���bØ��y�TO����Շ�'��e5ȡ��Y3,��ab��:5��Z[b�2ݚ�)�q?�"����5�X���|�H��e�y+�c���8�!��g��^ ݵ Ou`9'�����,��5#z�}�g�`���^ZM�>!� ���4�����Ƞ7������߾����l�i�l5I��
�C���9�S^�QNboa�8�߷�@q�xL,J���z[DQ��;��89�H�����Ş��ި�;#���dU&;�N�~�d$a�7��4] S�����.�  C�0�rF21�|���/��W#vw�*hq�[���$��<l���^6�>��:%�i.���aZ�%�Q�V������p3ὁ��b���7����I���oGߌ�� [2�s��q���Y��m�4��ߦܷ����ۊ�8�:0�_�K��m2�!]���W��:	�y( ����y�T�]w+�͡U1�S�M����ƜA�N��$��T���IWأ��iI��8㽨�G��.�.ԅ�h}5q��grU����9hF(���)@�q�a����N��>����-H��=zhc�؞,�44��[�g�T�>�Qp�|c(��T��7��]PP��#�~l��Ղx�++��1���ʏ��ii�����9m^��0�W&T�$SWC��pB0<�#���B��~	?'"Ҍ�w��'Υ@��|�h~G�LK�WB��(�_�Y��Z�9�=�L9�hGOn�7���M�����s�I��%7��s�t�����CA��;1}���֦��bD��`f�����4p�D�C�5��V,�N'�%A����M]����`�H���A@~߰l�"o��]�x\r��o��U�>;RORB�^��y�K}D])	w�YQ �A�s`��W�Kκǫ
(m�]Kh�3j'A�t<��m�q'��J�x�OE).%	$^R;!y��@X�=���R���(W�p�������!`z�슱���G��ɓ�@��Xn(�4V����y�o�
�&&���[�F+m��O�1q��5$U�|إo8���9���_���2����7B�#R����6O��?��� ȧ� #X�O1����'L�(rCH��c�G��V[3�����ǷeԺ