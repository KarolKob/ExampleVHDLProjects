XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%����]����7z,U������C4*Q[-����v�L����old+�z���$Pvq��������c�?��=�V-�*���q����&�)"��J�7��}��cP��=�F8m{���r�EuwbL0��73LnZ=ע�?ޛ���IK��=n=
0C�Qm�������φg�%@+��6���ĩҾ	{w���aC�}jNwႣ}d-���!���r��if�?�S�Ղ/������RtE��>ї�fB/.Zl��x�P���[0� ��Ŀ�3˨򦇹�,�ԟ�B�6�h�|�c�oW·*R�>}�26Kl豋ս���T�x��{	����רG���Ӥ�<��X��q4<ު'#u~���F�Z�GrpV�E�r�`���T�Rs��� �+�{q�K��kek粗�`X4WX9�}Jڪ��R�/�+J�VӞ6�lܢ��h��7d��:W�vX��I�jq�$LHn�2M�BV���[~_�����F�P�]?ǚw�F�2�y�	�?V�p;���|s�pl��Ё�\�3�D3���c�,l����3�g5���F^J~4�u�f�A��罊4T����*^N�* �`d�>�=��I{$֋���O��b	����OvS�1{5(�xʴ�,���Λ�����o�?^?�Y�O�;�n��@�8zE���`�pdC�З�X���!�"eI4
L��a��'�tK���|/T'���?<<6Wy����&ΐ��S�/��]`1d���=>�~��S�a��_+[�XlxVHYEB    10b5     410Ma�������q��`���� �-�g�Z!X>��ʓv�e�oßC��������Wű|�5>Fj�~����893�2��6λ;µ����W��Yd뿮�Y."p���f
�9��OP�wvLI.�Wt��24��!A��˚T�	��Zh9�qGb\ɂ`r���ˁjw$ �PjЋ���g��d�tŽ���TVT:�g`�s&������*Fm���}�,p�M�*ILx2��֎�at���|�.3z��@��v�nӅl��G���m�;�2���m���zm}D���E�3��+�EB������p#^�˷���>1�m�x\�.|7��zA6,Ey�L��D�2��ؼRt�T�K�$�es�x�x*�(?pQe�Q�e\z��7��Q~��2<���7w�H!Un��C��&��`2��6Q��E!�4进ş���2r�]�>�1t�^^q��h��t�9f�+%O(�M���d%���g+|����.QڋH��y
^��V�����U"[�<���c�0���#�r�Xr��:+���W=G$U2*?O�>O��0yV���Ç���,��s���q��e+���V�&f�s�&�gw(0�i�!���V���6^��tXu�pd�E�d��Z�C0�P��K$��5/7V����"����=Ք5�����@ m�RMS���l\��������cT[����Y^G޼C@���<���8��2��%�g M�s�*-[CÐ�'��@D�u��]u�m�o^��I�� ��e)9 _��f���I�^]@����"�090��)��qD��c���a���/\�rޡ;
��|�q¿���+����V�W�9�~( @�_!Y1��'2F���4�LqO�=;����ߨ)>)�f{��7�P��VRl:��R�K�����@��HQJ�}���Vx��<ˎ��})tH�,QJ�E���F�s��G�j�����,E�������2x7���mL�0�kؑ��4�z.�MP�_7~ٰg��2�Y�L��d