XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z�������a]�>��pq0����ѹ����9�@x����U�R���3��3]��`�� ��3���U��q�ְ��A�y���B~FVZ��1����z���(�z._����)֜�>�
KR���ڳW0�'�W�E,C���ZH<�ӊ��H��t;쥃,FAP��9�g&ު���侤�g2����_^��cٜ��Hȧg='h0��C�U$C/Mj�UZf]Kg`��Z��ے�Gٍ�2�~gͮ2���Ɗ�Z�-��
X�ѷ�����'E��?��d�y^�wb8r��v�G�ai�E�G��b�i#��8�Av�*��cS`:���M�V���΀1�]ˢ����x��	>櫈�^;�T0�	���Tj�Ң����L$c��s��/����KH��~c�W�����vo14��x���jIr�Ɵzb�+S��ӿ���� ��V'%��/W�.NNY�X��TD�_U�&��w�2
�=�"wǩ�H�&r�J��5xh���᠟��g�(��Lwd�o������5������D�2��b��L��#'�,/��A�N_���6�d�b��)ȥl�k6oW@D��;)�Q�=�6���XA.#�H�8�x�����s���4�Lz��������5�FS�zT�Dl��?����Lt8�i6#��QSB����6:G����kxV]2��=B�wkmz�w��Uۃ�����઼_���u����8CIe�V�-p�;o�NX�UB�V�tzXlxVHYEB     748     310��q�Ɔ��i*�L�i��a�^�Jz�X��P�zZ�AP�AT�L���
d	$�{,�?+B��'��������k��!���yĥ����7ė�:�d��16K�}�3��M=b�H�ߪ���Ͷ�g��b��ϼ%'�DS+� 8,c�HO�[����	6atƽd[�-�������G%�b�Jv�e�lsN�=�лcQT����"��?\X�$�i1M��f
h�P�*�,�wD ���g󅴠�[ܼ�j���,Y�bG�k-���1�$:#���p$�bB�:�1������T�����=�<�A�P޾j�Q�0�A�b�ͭ�\�wg���Ń���B.^>)�o[�{���N��{�w�-x�3~�"Z����Z�Ԉ�Wj,�a�&t{�ٰ_Mk�߶F�)s�?���������������%������A�P�sg�Tp�$�y"�?��f���弃����Q�Y�R±Qe�g�0_��*Lׄ]�%(�F;k{��X��z��ݟ=�`�2~��g�nJ���$y��wR��A2��mqup�;�1�#j�O���h�Cň9( ��I>�|�u��' �~�b��͕/_$#?f��
��<^��3b<�F�s�����9zZ������?�Q�I�웛����yB|�����>������#�(��p�(*}��s2�n%I|�9����~�#��~��	/��b
�r��KdҖ#^>��hz�O�^�%pW��¦���Yj�)���cMk��\�� ����GF�