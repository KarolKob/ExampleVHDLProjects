XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Y�8�>(�q�ԛĴ����7Aq?���Y�Ջ�E�3�pN�	E�M2"ߴAS�v�;��cS�����Te�B�W"�����NԎ~�� �)�2�ʰ��8�&�ء�Y��Uq]�t�b���PD�X��@Z4&��M��(Ƨ�6����B��pGQ�3��᭑/4b�_��F	X�K����w���~���y�9��9z8w�G,�B{L��(�����!��q�O*��Y3qLc7��Ԫ)�Q1�-��`
_Fr��O~��������s�"B0i`14i��l9a����G���7��:ֽ�^�{���f�1j��ӽe���*��OA���ܲ]��G��/�Z���<J���0�0#���[�5Y7:�n..V;l� �JA]�VgGJ�����h��K-M�U�q@w�%s����˼.}R؝爰��.���۞��Q��7ξ�ӥ�c����K94��T�֑7��4��Msz���(xP����N�xK����:�L?�]B\���"�N8�_%:*�|`�j ?�.�|Dv�yg:j
��`��]�)K��¤Y�S$:/ks̩O�������6�F��e#�dF���4�sFh���xO3�V�����ʭL�Y4)-��S������(�:Ӏ�7��˘|!����[7vk���#uj��(*�6%$}���<�=���k>x�0Q���Y@�L��0=\ǵ�]�iL�Jk�82#q _��Ť8@g�Z�Ǐ6�1DL4c7��XlxVHYEB     a7c     440;��q䆢q� 	]�+���:n'��Uғ�%��a�n�U�OPr��7���Mi8���I�����^������(H��)谫c�K���ha��Ŀ����1�$ ���훘5��
����q�%/���O��K�r5m���(?+U:�V��\5$���1r"�e��G���䵔��Q�u��q졣
�,�vb_����܀^o`�FO+�!����$82[A(�_�R��J`^p?���\��B���YZvV�˽ˌ�G<t�з���r��:�n�������"[�0� ��F����6wb�uD����ŭ����RY�������0�k�<�c�R����o�@!����.�bB1��F"��@�m���y'������wnU��*{~�I��u�t��P/:?�1+ɍ{�����3�>�bfT���,��3Ԯ1c֭8��	^F���jv�־���U����lK�[���i��/ ��T<�p ��mmљꉖ��l,N0��S�N�P�|�n��`*�âJ�>n�O�N�"h����av�ؗ'a/  y� ���U	��1��Xe�k���Ro,}4]���T��6"z�U�4T�� X�Η��t�m�6�܂#��dm������	ŀT&�#�2`>����N��q�t����e@&ׂ��HE=f�aw'�h?uH)f-�3=�\ǃaz�4=Os
[�p���䃆f���y�`C&������E����β���ށ��=q���H�UK�&�����u��il��1��-ϥb� �K���;�>�t_tnK}B�T"��__0q�E,��_��C�[	)-&`hڞ஼�4��2ƴRA��=릓k#�_��'b{�4�{C �fP@�R5�H�͉�/I�/TR�Rr���_q�zX(4@�˰-.��kڿ�T�a8������R�@^Έ��Ͻ�v~Z4#�Ģ�'�Hӽ>_c'Γ�����3�@���N��%%�g��VU��txl�p�@xl+��l�|�~To��DΘ*�=���>m�,�t�W3f�^9�/��4'��ed�@?���J�E*��I�}��>r