XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0gᖚ��tof��?~�J]��T�C��ݪ�5�|�tC�p{�X��K.�.�xlő��7E�NAs��+��#xI ��h�b��|wɛ�g��_S{���H����p�C�m=5��8��w&���eAą���'o-h`H��o�yG���]���&�ʹ.N�j��4������I�W%k���_�������#�+%X��LV����;��d���p�(ٍ�/�h�"��x��wDIHh����{G廯�o�t�|+�쮲#Y+������h���V� O�)��
y��nK��������8��e�)��PC�J<p�1~]�bŤ�n2Z k�@7}����̻���%P�0I�b�|/_�!���Edp�ڑ*I3�k��AFS k��c�0�wH�i'���UQ^��)#ֱ���mW��0���}mw��:b~^��O#(㴎�7��Epx�~L@���k��B��xE��a?�0k��f_y�Ȃ��)o��<0W�R��RPfx�
�P|:
�o��Pd,7}d�Z$h��SU
8����?�x���]�8�0���Ni�x*���=���#��}#W3�s�$����}kjFT�뼵YH�����9h��K#nk�����}��f!�b,h�n�����֛�A������� ��v�x0Nsd�u�V/���3��ʒ,at4lFA�*~�ʞΉ�Y�do 7)hv����w��@�|��F�-�DC�����XlxVHYEB     6c5     300E��Y�3������jA���GK�2���	��+:�H.�~~�+]'���qv�l�>f��DD���>k�e����ᮌ���WC�N40M�\���W�l��.�5r�9jmp�`�@�� G	w��v����3�Q؟��Z/�ӗ�\ӭ��+�B>�C9� �B�at����w�@��� 2F[g�����~��k;���>q�Z�6��S��^%gцB΄�>|�b�Ѫhj� R�ׁ[���4���Le���܀��+��'�l��*�c9Bb�t��ZH�uHcgZ�O�p��R�W,�"�`�+���¿`�ϗ���R\(�f���ߐ[�*}�u��ȗ��H/bB���3�%����c���H��P`=���h~�@B#;��[A�֪���uP�?��4.rɦɨ�w8!���V�W�-�y�<�QA%a�}��)ؼvIWC�%�?$Z9�}��,N��~��%C��]�����bYfYk���Lތ��VH�BL*���� �)�"�Nq�Ք���Qݭ���jJ2�j�GV(^cG��`���ZЖ�Z|CK������c���/�Y����O�Y3�@9YU�^1��-ݖ��U��9���P�!7���TМ);�W*׻f���C���Ք��M�<ՑN*\}�B|?&�Q{�&Z�C`=vE&H�<�	�
�Y�g�Q#X�%苻�?uHw�w`M����v j��F��!��x��#^�p��04� f(�H�c���,q���U�ǘ1J