XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`�8�������D����&��e�23�	���_������Q������pa���fPL(bp侶es�\
���?!���Z��|؝�F���Z��ȍ �����$���*S%��q�d�b�T�0��6��Q1��Ru�Z\�kY�	�.�HC��8/�N�ZU@�,�j��c�r�?�����ۑ}A����]��8O`�%a�L��� �eؿ�5�1��}�]�
i��u�͸F?��@j8�0��b^����d0��2�B�<� �agVD��G&0�~�8KS�-m:a��'o��^�kH�_��,�M�2��&]Y�c*S��f��4'ҫd�z��Ҝ��}��)�h���9��f&7U�T6�lt�3F�7�Ͼ�h�pgI�b04�ݶeGH����a-|:~�=��a�]����'�n���~���W2��(O��6/;#WD�'�b>@	���z�Z;����Di�k*��N~�c����b��yC4��T��>1����c�ݨ�)a�U�M"޹���^�jB�w�-$���B�]E�F��vG�K/�v��&�;>�r����ug7ߓ45-m�������8�)�28ٛy-_OU���p0(����$8���<|8A 3�̍�i?�":ҙ|������\��()��@�3�|��k8�)K�(@Y:�Ԣ⾂3vl�K}��R渕��λ��i���8�·�L�6����iŉIJ@�̌��5��R��2ӎ���sT�&U�ճL���r¢ژV��̮�y,�2� ��b��Ȣ�6XlxVHYEB    1621     410�u@��\7	�{�$�>l" ��O^SM=oKĩ���+�*ԛ|���|}X��O����.U��A��@q��v�Ѯ��P>���%�8C�Ki�H�3
�jN�9��]���L�f���,���3|�)�m�%㡘�|�К"nS��3$ B� ?�>Ѷ��4�[��\��Qk/� ��-N��#7fƷ�:��b٦�R
+O�~����-��sRP���B�2�#�&kTB`����%�hQ+
��#�"��h�M����؄oN�=���;rxW1�>'nE"�Y81��i�r����/Q��:�=�v�o�S�>Ԍ��3
�ţ�����>^��֎8/5f��#'b+��PXgNJ%�cA��kGb_e�㳱/�y�`5(��ń=g(�c�d���Qo��+slB�D���AQm��^f�_�S�E��]�x\�(AZD�9Pdn�|�A��T�[��b2}Vl���<���s�ݾ��`�D=�Q�1�-���:�D���/-N��5MP�X+]�ڬ�/�C��BЌV�z�S��U�T����M������<��Đ�DS�&"��K ��
D�)�`����idʧ�o�E�Ѣ�.�,_2��[�8�#��3���Β�Eru�f��v.K���m���$3�\�f�_L�tY_�h�5�ԯ3ݷ���J�	���*/�i���|3���v�V�-�(�A�~Q!&�`��py��x�������|m�*�����q�xy0�<�y�bG�TR�xN����;.��B�`�W%"���
aGk�<�"�E��|��<r��B��W�-��h����x.󏞪A��3&�c���U.�����H�?:��ֈM`���o[G�tXD&
��-�vm�[˾�}�_kG�����2�X+>r��Q��*� �M����ӫϾÑ�ĆL���\c�Ҷ.�2R�·R~���P2��'W�W�Sl�\���&|p�l�}p����@���xd�[ǫ�J���i	L�~,%��wB��o �cٙcT�U[N>�