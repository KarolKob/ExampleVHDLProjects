XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������c���W˖x\y�U�4��-cYɦ_m�]��:��R��D��Ȇ_<�M�9�:N`K6��g$@PN_+Z����rʧ������y�D��ҺB���#�������5IM��,DJ�#l@B*(��Y(��[xV��_���7��d��������xr�!A�8KJ�E�bݐM����'ns��P	��8�K�V��0.N��oD�UT|�25p�/^,��nD��T5�з��4��.�����"1߆/��툹��W8nq�)��^,>�c�4(�����A�U��Cu��S��Z�@M�)=ݺ���ڟ
a���a`���:}4̧������e<tƂ��@W�2�9��%��.XS!Y�xȾ�S�#�P��P�˔�~,I��V��逮&����H���,���Ϲj�������
�}g#�I�%y{�Z�H��رsWA���B��}���=(�'��2��U�an\e?e���0"�v�zR<��[�erpO���[Ic\�w$Se���K�Re�&��u�^� �%�k4S@�*�R���>CS|Oڑ3����! ?���u]���[h��V��H����
����<����놗��怃K��4o~.�8��3������ə��E�H�P{��AUo�µ.�L�#x4$s�Ii���:�D!|jk�d�jK[��So.����a��PRlR��<�CK�o��$�0��M�7D���n}5��֟W�x ���Nbj�B��������2KBq�XlxVHYEB     99f     360̨�&a�f������rf�{��2���nk{,\��z�����g	M#�$}|�Ea�~��b���[1�D�`F���"�ڜm�o�Y���@�ݣ��KC�:}gr��O���<�m�ؐ0������Uƹ���J�{|N��`�AWo��7�&�Q���J`H����'kZL)S��/#ٲ<�{Wl���)�6�z �̯kϺ��A���¼xU��tZ�}qkZ�}��f�k��5!#���V��Z[R�0�`���J�~?�s�L��a3�E�<��U.ޮSo��
�'ߘ�!˵���TZ����$^�M���4Q˄�P��h��^�V�e��?� ��a�ĨPO+7�n��Xr�6��67�\�SXo�g�Vћ�t/�΍�Շ�U�J/�?��Z� [�u�s��v�a����Y��}UC2y[������t������z'��]3ZQ��\�Kk�$�T�8���0eE�MV��8���TC.����wX�ѱ��G�-���W1�O�FxK���e
0Yg�M��7Ј=^dl6�J�������֖��ݤ�ũ��u�t�M^�F*ܴn�4:޼^0/��,5���ZA��GmZ+`���G7H5dvO��S&����"/ TX����WA�}���Vq2��,w��X��6�4�p)*�E5��N�p����@�� �G�a)�a3������.ۆ����@E���`ѿ��m�'s��i&��Ym�7�4����K��U� ,`���[H�c�Tn��@/S���s���@�E�|����T����u����#�{�i3qR?��~��'ـ#+�'�:���2����z��E�+�rڠ.R�=�	��c;S+�Zׂu�b]