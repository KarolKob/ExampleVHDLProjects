XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:Z�Ss�l�ۯ��B};���K9�^��ĀG;ee����Nӆ?���zY&�ؾ�aYVX���1��f��Z�+��r�P���5�%إVh�I��7��í��L��{����a�擭\7cWg)-�G�t��U�]�Ğ~�+���B��ĒmQ7JH�4ت�C�/o�|���-�BPG��ncn�9�����=偼�T���拓E�.Θ��K�2W7ĘE�z�\�����E.W��mCCݰ�ra]�6���Hz7�:�ʃ�T��x�k���� Q&�qQ��������O��C����� V �p��f�f�ER��/��5��G0e�b#'�9�Ɋ������F+���';8.�E�����d����w�J��f���ҷ�w5���·����5��Z�7ڠ�F�����F1x�";7��㟉h[ ����n%�t���k�N�z���H[j���sr��`��_�Γ�#B������r2=�������p�4mޣO��p�2��Xhx�e�a*]�Ek-x�7��N5����]�^�
f݆�TG�y<k�Ɛ���y7H*m����*c���桎Tmw��<@
�/�8��$�����g\�ڠ�M2O�NQٍ�PX�H����TmˏQ����z�-/�e��7s��
nuݝV&p="#߭���1�i���O,j䌣ރG�	�� _�ĺ^N#ˢ�8۽3R��W�����t^Z���"J=�W�,��NDh�m:u�O/���"(��a�,XlxVHYEB    60e7     cd0>�7����Y�Cka���Ƒ^7X&�E����Z;`��?���p�� ��(���%�H ѝFۑ��{#�Ql66����.��^��J�J�q��I�7I��S!ݍ&rg�g����X���I2R�,̂V*��tWP��o��EKb�w����rq@�i�b��=��T`-a2'm[�+\��r�t)U���gU�.�{^��]|kF\��@NMtr[��I!wv�%�k��~����SMϾp]�/��XCn,�>���� Y�$��v	�(_�n���S�O��[��������K:��.mE�5�Q�����$����]D2�g�gt�Xe4��H�����+-�{$�r.�(
	 M&�GQ�]����r,�U6k��T��1��)=�䬾u~w�$�7y�!�E�0���и��W�!R�Tt��	��e���%y��]<
�&��˩gS'څ�A\���&�久�"�"�hqNo���6G�ѠY�1�!�K�Zv�U���x��^�B��(5걓s%8�{��Z�SJY
�u�1�U<�W��4���v��e�bVlb�Ğdc*ޚ!��f$R ������p��0�@��X����]�0f5�3�F���r�u^����g'Q��xaW)����D4��=������Qp� H���첋 ���¶�n�,(�(�j�FC��%΀V�2�0H��Bʮ�j�{���ϖ�n]%�H��#��(�ʑ��Fp�wS��gc��1�����V	=[�ɞG�)�`����9��I���7ɸ?�Wa��B:H����-v&z�l��z;�]q����JE���J�a_W6�#��k}�4�����M^8���@��2^%�m���Ӌe���"�9x��A��ۯ~}i>���@FT��à��T\�~�uzט�5�\��q�@ .ޞ�^N��\�I5Z�+� �0gd*跊~E�5	��%>)4B����}����5���G�+qC�3���G���Z5��b&�H{8'G�M`y�{*�-���V"af���C!jp������-�����`!��:�u��L��A�01^��O�+ ,�[k���aUX00��,慡vs��?� ,�bydɍ��	p��̷����Y��)����=޸���3\�Pq��eje�露�t��xp��"9��#�u�ƌV-xa��P02/�M(EY��'��Tqu{��%����,�Z��|�a).N�󿮦y���`c�,���K�����.% �ktjO�̈>��Xr<��
�����ՠ��jg���PG&u�^i�] m���R�Y���w��`k�������l�px����O��?�P#�?�V��:���K�{z#�]҃���D�`>�N�we����+����OA�ݻ�㸫@q�
�dc�y�J0�I<�G��Re/Lj�Iis%�?�E � �ă�[��$ w�7���h����kF����Boƥ�^*�z����_�ZT���wWY��)�J�	s�6ʧ�0%��R�U)�D'/$�o�u��|'�}"ag؄ڀAu�P7rU#&<^��Is<�����¬���4!����r6O�޹�=���W5������p�������M4r��Dm���u\�������`T�Kg���f�Z RV]ǳ�a�N�	m�t ヴu��{!|K�\���}�g�/r	
s�	K��³,�%e�1�%ڤy�B����6��]�֭�M���f&�>z�)[��l`�NZ���]���:B��H�#����g ��,�� ��̹��
�����m��R�˸2���fES�ڳ[%����1(y��{�t�٨{��|��lL��'��D�%N�>�B�c���S!��y蝵��;'��;����gR&+C]ms�$�HyZr-�ͤ)q��nG5�P*�	�x�8*f�����b�Z�ԧ��ڔ2^��uC��T�mw��,�yv�n�������F5����i�DO|�A��ͧzv��BXAc��+R�t�0�º�y
&�5)�b*�]D���fro-���>;2��[\]����\G�;$w��K͍�!�7�r~wa��ó���/�Lݫنd���A.:��Y��-�
}	�6_��Ӥ�"W���r����?ގߡ�ҧ4����<iD��-Tf�DV Ɏ��P=)n]y�,�t%�E.�9�ˉ$���2�������ea2S�WU����9�/Hʋ���������j�G`u�z�NW�N�u�
���'��	���)¶
$�	~��`r��1����%�۴��<���E����D6X|��~�������TFsyr�U���͍1R���e,ZJ؄��V���Ga�u(J��F�DO���J�Rı�q�9���8�66M��tK1#�^t�8;V�� c���C�j�UE�������-�5�0�;�)�+p5�3�=^������M!gT9�|s� N�����)��[S��a�js��˞_u�es��T�we{����N��|2=���P;�)m�ZU�:/�ւ�Q��+g����J~�=�#+������ %�btu.���@w��<���q�L�"���})��~/7�E���E��h%� ݖƈ�˛��bI����*>����q�ak"�� �ۓ�Po1��w�-|�� {p�fE�уj�3pU�%�"�?�e��Qv[�I;@�{���^���n�0�ཥa�#�GNbky������MH�!b-�*��mE�e�e�_a��/4�{z����Dw����Jt�@���Q�r�Hi����!C4�DQ{'�z�E����|ާ�,�	��IW��`�n��i��}�XC���G�0�x�j>�u<Y���n�kP��n���jϐD�iK��H�t�M���΃�6ف{��N	5l5��6�DC��w#�Q�9V(���$���1WS�S�vmc_p"���+[�#��+02�XΔҤm��c^*w}GQ�XT6[q�Tg���&��s���Bm�@%�Q�����)�Ǵ�X�1��6�4tRa��u|�
5��T���.u9jٹr�ib�ykUsM�z���R�^?�w'�������6'\�EOt#XV@Q����R_����Trj�iV��)]�ĉЍ�K���I���S]sc|�����E�+Ӈh8��%o{����=�[�ĕ�
U ��
�Q���|J��{(�U�ʷ�Y�mu
�uSℰ�Ϋ�ϖK.�YIlDX����-�N:�w���,ɂD�+cY���x|N_�D�xs��	�Ɨ@�5��	����bL�{}���A