XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����PQG�����;��o%e���c�h(�W�C�q�zu*S����{p�2sza��q�Õ �l�*�7F`��0r��}A�77��W�i�p�Ό�&Dcq%I�}��%�/�k�P`q���� ��G���{�?����i�˿���4�P{Ch�w��q!��"�x	B ��ynU���<����8M����M��y6r�H�m��/��;�[ `����]-	���! ^2�n�u�e���D��[���)$�W��Z���-'X��%I -h�D�:��t��w"��s=)���P�dh�h%N�^E�]�HC�Zj�J�xI��%ف5n�Q��\r�nTo�h?����D��PB��(�0�;j�� ������Sـ>{��M� %}��4��1�%����AS��x8\�GJB�q^���� �p����6;����>>�ā�A���!#��^ш���F���4�ۯ�������͚�܍y��\�Ĩ�\ڤr��DWz����ϧ�V�*恤t��=%����|"C�D�q�Jk�&b�cQrI���-i��>ı]?��`�l�:��_�
��-��r�nM���>��&�gEW�d�V��h��	8~Hݛ;�c0y�G*�G{|�� $�]�D|tA@��"1/$��_3��� S�T,�1�z�&�p��+���Oj��	Q������N�:��\[tEIT��I��/S��#L����M�5��V	�{�����*%_��k\��J��v�B�f$ǚ�F^�XlxVHYEB     e3f     440�_c�f<o�����E�s�����m�s���	 �x	�ö�8XכLI�_�'XS��{o�-B���@�DO��Ȯ&L�Yb�p��+��W�j�a=B�m&���M�m�wg��PِQ��tv'T���Z=y��ö�v�T�5�Mk��3um��5�^q��_���C�8.��]�
:�2�M�W�#^R��T��6D��@%?xH�����o��Ked8�w��~�h����D#�g]	�j}��ahQi���P,s72u%�8��X���Q;�M�5��7̈́�r:@u�5+33��&�ߋ�dh�HBr!vq@DP�ᄈ�b�H�",�?�K��㙸IJX�P�uUn�n�Z�۾So!�'H���-��A��hZ�?ք$�J�5jQN��C�����k�jȖ����M�-q�-�EZ���$�]ٙ����dj�;$�����v�7�d���%[��� q�����m�n]�Rڼ�U�>	֌����D��Gx!��O1�����T; ��̳_.�$|u�vfF���$zEV_�[�X@-�N�E۪r��Aq�T�~;�a:ʎ�nL�Y5�����G���a�y�8��_��FЌ��4Þ���0XW�[��L\�+�f��}�PwH�Ξ�W�'��b1o����v>9�!a��*�̿����ۢK�V�Q�c���
�4m�s�B��Bھyv�p�]�=ʵ���ULŭ��žRbV�fN`�I U{s2�UZ�4��'
,9Th`��Ж���9O&��3�Ǻk�U�d��^�@k��)�"��d_
:�`�i__gt�ԧ��x $��TR��\�Y�����a��k5�P{��Q�F�0h�L�\2d@T�H�Ô�	A�P�[Y9��]k�K.{��ץnJ�GŮF3��/��.������yu�W��	]��Y)$�$NKy/b��m�\m�t�Y*11�l�Иռ[%bG�o�k��>
����`�+o�,f#�	u�Hpҹz�i�%A������!BܧPU�K��Mc��џw%N���e�TE|�7�gS�x7ftIx�ud�{"W�*�缨*��t���燵<S"*