XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��MS��^�l+�� ���O���WQ��ta_���E����JX�)=d�s�M���^�[;�"�e�W���S���`�`^���S<�d�\�(h�����a�F���\�^��k���TB=��R,���ݪ� ��NQ@"���,�֮Hc�_d��I�/!6<;8԰�
�-f���>z��TY�N�ʶ\���H?3RPIpq���@t�lx�q���V����r32F��9�]G��d?Д�q���r�QVp3�k/��m���=`|
�S�Ykև�/Ԯ!L4����I�۰b�HS�v���3_	�	X�$�݀�~�ŗ+x:e2T�pLg*��ȯI�q�m�Ϧ��{�%�L��}��gP����#n��h��%!����s_�u:�2xm�O��0�㻱\�{֓�odU�м�������r�Ut`����d�ֺ��:kr�t��������ծ��]�`�����u��9�Ngoe�6TN��]�[��Y����ո�xӐ�xˎiN����&巊y�n��{`�!'A$��h�fcFO�"���!M�x�e��ɦmL*�o+���J��Xz?��h�ģ�;'MX��/.��o�P+b�DwQ@���]x��g�jo�f���uy���b�Ȏ.�0���P1��C���oP\X�\�������tm�� ��Ë6�����N��Ι:�`��z���3-��;U*#�����a�ۃЗam5h�����}�1grT���c8��ŭ��XlxVHYEB     686     2f0u��e���Bi�+��/�#�ky�VHo`%PU�	-2��'�{���6�R�3'5M\*Z�:�4n9�\��ZWX@����x� �3R$�lߋ��sJ�\�B������e�O��F�����Y��VP�60jMf��T�5�D����B@(r���H�Z��1<Gw��4��U4J��7��7l0u �Q߿�����v(*��b�����j7Ďd��v<{���9��-�Ϝէ��,X����~���޹	���JB��b�^Ն�Ƨ�f�d<t�HK�Ʋ��}L��q(Ē�X��CQ�8֡��[�o��ɳ��?I"����f����S1�@�o�Hbi�����g���*5���"�0����y�������
�z�K���tي�}���G���4(�a���h��v�����j_�wj��M�e|K��B��̼�eΐ��^�fR�ziȑ'U[��i�C�Uz6��|1�Iǋ������U0-\�(�U���x2 ��� �|�7��y�ĢL��E5td"h;Rp��K�Z͡��p
�A�V�>|F���dJ�Y�8�_U�@�(���Y�)���Ʈ_�>�vf_�>̍ f���	N�`�`KU�}&Fq�\9H�0�$5)
�Ɖ.ζ�G)+D�@��S�z�î.����P���2:,�	�&"�:@5k<�2�H���#��{���E=�Ґnn��l����t��� L�v&��k�8<�)Jp����88���Y