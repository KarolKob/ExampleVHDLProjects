XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����� ��J���̰��Y�����}�~&i�y�����c!i)!�;oc�����[6�~���\oRn���=N��IT�Rl��m��gu!�83ii��1Ybj
?�F2#���c�+����E�-�Μ�P���pD��I�zi��[��b���2TLT�ϔV�x&H�y_ �xpsq;nrݰ����cI=ڰ�,P��[�H�����Ֆ�)e�X�9��کs��!ߨ-	���Lε��+����ј��o���xO� 8jf�,%]HbH]�eP����Ojo�{�T<[Rn#���(�!`80�R��><�Nd�&Ōw��Ķ@T�Rը�J,��(V�?�3S�k,D~�j�*��3w�̻���S�0���6�M1>����������(�G]��6�S❿A�{GO�kt�����oIQ�ż��c�s!7j�?�7@o�r�slXr�>���4�̤x�bmc�Lm�����S�s(���/%��6q8�;!c�O��~�r�*�ݙI:k�,�1;��H����*�!/�A.'x��� ��K����Iȝļ���+:�UD�o�7X��}W:B����A˗	og� "NG���?|6ތ8��|M��j�8���w����x��J�N�1�Sq����,�v���IZh�������F+k��2�� n`��bD�M_���fe�q�� ��R���wk=�Hs�dΗ	��Dp_׏�χ,��`�LW��=��a1:�q�d�)�BE���XlxVHYEB     935     3e0�%R#���t��z����A��yӍ�#6r��fR�p���jI �XP��9�j"]��tkdí~HԏUcڹ���Ėem�`��9���hk���H�!����?n�����d�����WS_���8���xDlh%7�v�,��;�Q(�-�4��s(��%Q�(�Hm�n�{_5��0#\ٓw��-M	��/@Ӓ���RPf0p#�C�?.�K�|�-P�`;B^a�H"1Z���Оg�dA-\1BJ_�̻�z����'{ߊ��wno߅[�e��e��hL��X�����k�H�^[q��O�N��-��Q�E�:�y��wH�^��=���b�2Pu�-_���ܟ��_'Hѐ�n���b^o�N���Qgڦ��ü�Oc9`,.�}�MA�ב���@���g�,��|���&N>�f�;��2 _��vM�"l��F� :;��<@�qJu��B�eT��B%9�{	�=S�#��!��Xs���Z�a�Z��b3��L�5#H� ���hǥ�洓΂T�rt
vT�P/+���s�V���3`:���(��*��ۡRȕl�7$�YE�H�?*M}�o� ��B̹3K�@����Ja�ȋ�0���'ἂ�DT����ZQEu�Sf���;��n�
�x�F�w���fp�����'m=ȑt�k/r�}�e1	1�nK13x�������[MÈ��n!�e�턜Q�< `�e+5�J4^k��F��ځ�m{�7%�K ��Zl=?�W
s�}ZU�{�.���H_�,O��J�.����V~������/fN/a��	ת��=a�xs�S�����*�Yg��gT�2���I �P����,SbP	����§RE�y?�ϡ�����F%�,�7��.�GO���'�$�̠ȽU˭GY�h�ݖ�|˿�O۟�[R`}����*��/�i�G��D���J�+�������7�qy\Ά�����zq���el