XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����,��	�	�`i;���B��;p�Xț(�]J>A�c�� &A�`B�����(�զ��/#�g�������S����J!&����K~j}�)bO�5s%�.�G.#��ѭE��Gc�6�n����8������qJ2��o	���E�Z�m��q3�鋄��&�O��F��G<�K�����B�^ұg� �0�Ϗ����H���!�{�W2� �2�>��D�s�����!��I����ú"��\2��_n�F��0a{�vrz�Cv?�v�9�z��FA��A1]}q��H�H+n�%��lZ��VJ>���|�E�EP#�V�}�)¨,������x<�5jx�>K��og3�T�
9tW�yQ!Qd�e%U��S����@/n y̸��!M�#�I�:�vo�k�e��2�Je��&�csi���*. �,sX��E��W���s�I�����x��e�K<B¹.�G�]�ʩ��� -�����Yl�Ķ��*���� Vn�4�!��筼P՟�FiӁe��⪋X�l�`�[l��b�W
%=���4cG�۞����.t��^���>��y �C��~\�߂���W:DMO����]��`z�a�č�l}��j���>�����HHI�W"�|�Kq-S���fB�XuW+�;M�vE[X"��%�ҸR�[�K��]
4pq'*,��&�I��Y��9c���� '�}���$��й��}��|'s[MK�܂&s;�0�l� �XX>�XlxVHYEB    1d56     780�h �����<�`�K���,݌��N�n[y�x���K{d�hH��}�(�8|����y�������}��^M/�����Y��əą4�;mǉ��Ari~��`O������別��a����'Z��d|h������¸��9w@C���w��bz������a"��T�/�����q�H��93\p`?a�(G݌);^_Ud�c�gk42�|�x	���/��1�@� ]��|���n�>V,�
�DS/ҵ8o��,�c�y��Ő�i�4BLLuA�4�K�C�_�U��a�G5�_?�S����Bk�`�G9m
�&}�lSr�4��a�K�����6E�^�A�'5t�z!'4��	"��$�hvg�8��8�`\���*S�%�	B�A��,d�
l2��F�j�|m�N夤�|~b~Ud[��}?�6ULِ��Oj!�e��$��<`��!
)V���:���nhD']�sE����ȅ�Y�.�}E�^\�%��ܱ���%M��m2~-�d���%���R!����`%��,ߎ��K�H`g�]m����$D>xZ<��:&��zEH'���u �z	ʒ�����yv�lﺰ�{��.Ezo�=�N�N��̹���z4D�-��z`�¢�r[�@�&?���������`�@o��k������L����1���ejy��n,��.%���θ�ŏ�z�Ar�����S���e�{���!��O���Ћ��ނ�m_h$�_u�5��|����K���/�ȏ��U���z�ݕ����z:���1�3��ܞp���g��k7'�oysr��@Q����Mv&����}鮓��,fb#hܢ��'�*5A�	e(di�u��.��ӆ�b����Wu��u���'��,���K�?E�����M�.G��E��\�z���{��▸$�h�����2�-�1�9�R��rh�����"��ܲ^���Y���4.L�v�Ci�����/�C����w�����ï�n�S�u���؆_W��4d����'b!�xy9O��/��{�"�=?�`����k���E�YX-��XZ�r1� T��ϟ8��h����~�r�C�Z2�td�?�V1����,�V]m�����3|�h��I�Ĭ�`B2fi��حߙ¸�G̶/�.�XU㴍n=m�}�o�I�N�� ���[��$$�ł
�����|�k$(��Պ��+s���g�E_]dY�p�s�aʁFJJEdkb`��$z=M>����:>����w��VG�I¹j#9ջ��&R�%$+[�N��y2�oIWG=��=�v̢bܓ~h/	dڵu?�z��A���Oi�{�@�G�� x��la,�S\G�<��/���3�4��dS���</����N��Ċ2����` .�2�����%<V3i^�X�S^̔Z؈�8$Gv/�j�_�A����30�슿�K���S���#���K�������tZe*��Z*���1���UjK�-h,ۀ��$r�"=���_}ՌMS�J�G�@}Q��H.ۄ�J(���hw-�N2?օ~6�HI�Ʉo��@��?KG�L;i��C� QM����!��[�ȴj�˦i9k9�r~B���͖Dg4q��Oa*&�=$���y~�5+�Qg��o�q��n,�Z	�i�j�5Ds���r�e�{uO�9cL�E^̖��j����w���@����r6�|@
v@0����n� ������Uz��{���Ix9H��0� �2p���5�cF���Nj�!l[�:�6�	P�٦%B�fr�5=�<�L-]F��_�����y�$3)�o��W������a^W��l4�k�!o�M�T�����/����y,�^��^ݠ,���Gx����|��