XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������kLfN��~��;*rbʪT+�?���b2���$�F(��a�`���C���/�%V�Ų�4Rgy�fz����F(�R=�������>;\{�Aw���W��8��I'��á��U� ��º��"EJ'�aNϣ!}y"��՝Q� `��'mñ����6�$��jB�7I���w�_Wp�6�s�ȡ�-���n���q���a�HH�Q������$X�ly��. <� ��?��ɬ�~?�n�B�Q��?�i)��/��_*N�LT����ޱyӻ����Y c:/g�r���%ª�p�|Ć$�Ӓ�k�:���U1�ԅGo�t=b��z셰v['�T��\��̕iͭ�݌mߨ���s�'�C���i�'.N�O�8��tn�~�C�w�i�9��Ywm��V�M;.��>���S�ܝ[�F��4�V~�U��Ï�q'���!QU��{KIU\ؑ&7�/�;/U��U@R��I��W�;x�6��?��S�W���`v�S��|k�[����/�^Y%��|@�M�)��݁�鱋+΅���v���Y�3�*e$3�RŒzG�<���9BpR�!a�W�<��z:�7
�l�NT��HZ����v5�*�M��]LAy�ۗ�V{�������چ� 	x�������
��"Rݓ�Z����)$�������ā��9� y;K,�K3hc��~ἳ�۴�o"���5�&瘰w� Q���!oØ�ɯ>E�a�Uƽʮl��-��T��)�t����XlxVHYEB     b8b     3b0=���ȩ�M2�ZjjY�NHxD�����<7�6��[�8.D���ϧ�C�1�_�%y����!�ZTM�E\���^)o�E�mWV5 �To��A]tS�&�
��������E��¡���w(U���UU�B|�@��� �mSX�8�j4`%�ۓEx,��i.�_��TX^��%�8��S���X
�9מ���nŞ���<wIW^�k�kcG��.��9w�� �0�s����\�z��m�ۿѽ������7%��W�p`1���!��2��f��(6�g0GǢ��Q$4.��7^7�*��bP���8��������W3��
W�i��W=S�9��X v�Y,���,��,�x�<f�0!�U� ;�����a�����6�L#��6D���!�*tᾡ�
񗱔����%$(X`�ȋ�B}������ձ���^'%�v=��cY��[1�=*x���hB�5R����D��!�H��I���'
��zדt�?i��j��Y`�d�[�^�2Wΰ��*@����~�ּ{����+�3xf���<1��i%vo���.':�C�f��?$w5 �gX\��5�O�?���fH���"��FFu�V^wv��;/�z�}C�{�Mdq=#���ݎK����7�e��z��D�F�+F�����d#��۷���KG��)IěO�Xi��|c�P��.gv��Ir��"�;�wN�ǒ�!�����i��7�3�ײō���!����[Ĩ思�3Ӥ
��m�2B*��A�z�]�{�^�K��#
h`�pv�4(ef��N}����pW߭d~�L��Ya�^�ج��0�����*�@��6��e�5���/k��y�$�@s`��F����Û��Y���E���R՚=5p����l��#64|�P"K��ˡ1�s��WM���