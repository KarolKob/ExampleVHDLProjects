XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�oQ��Z��U'ހ��V�xp$s�|N�3��Ƀ�2(���v��Y��]ڮ�m�J����(�����H���s��%�>��3��+�,n�t�-���{�o������u�tp�0*�L*|׌`��cׂ(���ж�S�ɞ��Pu6C�Xw�����_����X<k����ڃh��w+?��������D�a��Ƞj9���a���H��>[�Û�͹e�z�6qNHj�d�,�Lߪ�/��Ѹ�>�@R��|��-�m�S[7��FG�A_Dq^��@I~���<��&�V����E�Ĵ����&/R���u��&�;՝��"�)9�B�H�c	G#�z1�WaP������s��t�&�V�y�����%�)vT�$n�z��nP뙿'ωEB)���kX��"sg't�!n!�6Q>���Y^�h>$b�.<P闸"�������Fy��L(�0�	��8.#|5�_YN{�ӓz5}>O�]�^� O��W;PQviB���h���&��|(�,���1DP�
��?����Nmܭ:>L��l�ҟ���:�KDXE�������4���z��z:J4��Z��d���Z��3���^�-�q$������o<��=�<^�|�hba��9�='xF����wZG��u?iz��&��N�#�I�{��������x�/"�f�=�f����qI8َ�)�X<}@�d��X��p؉@Y�|5��H��.UU�n�e����XlxVHYEB    249f     6e0����wMnN��?ao��Fߍ�pZh�Ǜ%
��kj�`�@"�to*�"�8����Ft�2w���D�� ����/T?�
`+��L�D!q�\/&�B�;�����7NH�}�b��e~ O�Gqjr�K)]�+�S�7^N]�^�Y��"AK<Jx�4ڼF"�"��a#�KN���Fy�bx�!g�e�ew�S�t#/��_5F��C��-���D����lz�4�����;��
.�K!����R��'m��~ad�x�N�g���3v��#>��P�Y��=����J�¬��D.��J��_�r�Y����??�f���7���ޕ�U��U#pM�7-:"�/g�ix�(b��q%R�>�R�^,�޾f�~`3G �	�^<Gsdp�����^�F�74�����*ힵW'�Ԕ7)?�K���1�M b���Jt�w4#{�����b[z��Q����ƌ������k���Rvr�uq
�Vx'��9�M��J9�!US�2�o*L߾���?]O��
JC>�U:̨�1�E7��PZ�쟡�dÌS-�u���b{�'7.��c�~�{���5�a��6�*����;����^�c��a�󎐯�F�����ġ���\�s��B�r�@���z��m��&�Ӑ7MS|��b��|��&�-������T�Lf���;߳tδ�-%I�xe7�3�����
�7aO��$����]=��?ٶ �N{��ɮp�4Dk���T��:a�W�e��&��S��[9��؋XOQb��8�(������f��}
��ގ��w`y�2&�:�6����m���:Ϩ�j�XZvP�>��)����O2<jEP�p˛�L\Xl��Zc(=¼�9���,�Lh�$g"(U\���+3����1�Ebb�m�?��G�	����@>�˴� 8�hb;kg�hH��ά[�ኚk�5O�U2ۄ��tĸBE��ց���ߵV��0?D�*�P�}[s�\����N�6��b���"L	}�2�;�{{���<^վ����@h��h�F���Ҡ`����,F�O�|6�`ֲ�������� ��U<�0��>Z�Z���$��[���]��j�)I/x4�d�Ann�B�ğ��y�0=�S'I��Q�=�=Nʔ�G��L=vXn��Jz�D �?0��H�x��n��{��9(!��v��gL��k��⮴`�gPx��䚺z��NK��iPp���_M>�7	� �t�Vp�w	��Р1�vd4Դ�F��� ��(5�nEVE,�>�E+�_ʍ.̩���E���.�q
9����E��:�G��R�Aԭs	��E�8$f�R��a�,�=)P"��پ�R��b9D�9i�?���P�U�m���}�3�*�\a3θ���w��oEi�iJ�r>+;}�8e|��5�~!^����j]���v_�?'�?]� ��Inu�+�?]�.:i���:`B���̆�0�)C�C��.TgZYݸ=�Ut�c���ςp���P�U%��k_�P_B�{�jY}Ѡk#nG�*�D��X�Y���ܷ�U:��6��ͬ�J5q�΋�m����-!�*��D���h>G�0�cx�V�;F�D����K'_1���źd	�}�e�Y��1r��e�W���kU��#_��UD��9�o��4��.��7����_	1��>H~x#��pTO��ͧ����d8<T�N�-��:ݖ{�}A�UxO��.�:�[+�����>�//�)jo�@���8-�