XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������nY[d���d��o7.���qL�o�ov���a��'S�i�~Y�h�&Ê��zO��U����J��
ʀh�SURq��ʞ��c�\�ם��L�k��.��Y]�Q�c����.�5����
z���#/ԡ�Hx'{LfIV����=r�Y��W����{�ԍ���#�M�L��[�k�^�ȸ��֍'�EM_��$2I����Km�Xi 8�6�K*[�=�^��E*!�ê����9�KV�j�� �&<�l�k̖=��:c|B��m��2����%������L��f�P`u��-Ai`o��*#������ʳ`>(�e��sV���8��(�C������0�+$��ޢ�m|�A�&����{���!8C_V�2˥���{.�a�V�� ƫ���+@�26Y�͏��U��8 *��p�I�bXk���Y*K_�>y���8`sVn��
����'N�J�Z ��̾��c$�8{D8�S*�w�������4e�W@�R��B����S��O
��&��=<�����3���A�h��A���52f��*N��\M�ՠ��[�(� ��?�������EK�Y��ܵ��0�o�U+HJ��i������$U��d&�r&h�#�o�y�*������E
G/M�1���1�?�����H�cLf�C����:f1*��9A���)�:�$v^6V��oѝ�ⷳ�φ�m7����~������v^�3M�κ?����������/�����b��멼XlxVHYEB    1c48     560jLh�P�<Z+�4�?YC�9�wP���J7���B�Q07R��P�N�`��o#����{��Ǣ�q(�"�Cw\���g~�&b����ҿ��Xhm���V���tٿ �P?�6h�RT���`%���'�F�_+��F�բ�S`�	r.�+T�J����c���.�`!Nv�վۓ�nٕ�����P~Qݒ�6e���7'b���\Ly���v2)D�jm�՗.�u���U��̭y�ngg�I��T`�s_��*�(S����-ȣs�E�JLr@�;�s��/��N�Ө���!�5��n
���3��G���>G�-��&'`��h�:P�����E�ݾ��f����]A��4+&���?R��~Y�}�v�I���x$;)�w�񜷝����$s�rp�?i��<���dn�=׼c�i$|�(P��hρ�U�S�vJ��d�R�7����}�H�B,��ͤYl�ј�.�'��q��_h��q���`�$#�d �r�f���-1����;7v��с"��<>�;��>"L>��������E���ؗ��ʍ�#�
q�H*�Z_�(���?�61<�-�������|��v���E]>��/�hdF׫�	�L�l	�MX(��]hn���5�Z�?:�)�Àf�Y��oDS�/O;�F�c܃���A@��M���h&Ml�����	�����P��M6�nR�>��7z?��~>&�:"�$C�_��Ly�#������j���RW(��Qv ����ʠU���!��Y
-�c	^'�bw���\k������|�Q�B����y�ȁ88_]=�X?#��4�xN<���$�M	�(*5�b�müٶ�I"^�+�p-�U+���I�O�d���º�*���{D�A���m�h7Q��d,���:��?����VW
{��ȴ���(� �������*cj�/�a`�
���&c������M�GZԄq��Yϙڐ�˒�Ƌ$�9��������LM��2�
i�fVW�F2�&��5¦��-�c4��o#$� �Dt1�����f�����kN T]S�p ^{�5�wkGB��I�\��kK�6�q�]��_ �L��Pe�ПH�$�?_�l�������9��ꪘH<`��?�e-D��cǺ���o,�9�<�f>�N�G�f~�R;���S�������3������|���v��7*��_���<uJ+�Ѻ�e�Q�"�ȩd��[U>J̷I0�i�=-D ͏{�@�m��z��+�]�F$(��Z���:����ԉC��'S>`��u�ȗ�lIN�g�h���4�fk�T�䓫��oކ�PB��`'c�;�?��I