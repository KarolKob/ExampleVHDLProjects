XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ao�QN�>נ�\~�z�u.�Q�V~�kQ��f�^T���ӊ�.0����I6�|	��{=�a���t����yVM
˻!�8HCdR��=���
���.��aL0Aۅ�q6
e�j��|��1+���$� l�%B�ӊCU��U}�)�M��9��=}~����g��ra�c�.�T��� �)a���0�t��7���=6�,���Lګ�	hg�����h0u}�	7�'������\�M� "��j�
W��ud�s�A
?��[I\�"?�ug����?a7������}�0�o��/&�)-���<�j���>Rj���i4L��T�$?e�M=s���X=�TU����|/��n��卢n}^S��n��pw�GSߪ3�8�5_��]�r�]�qi�'���0����B!XC�o�c�(3�vv�'1�T�}~g+h��,���PC��^��V�]r��������i��^�b��Swg�l����|]�i(Ǡ*+wy8�X˘�l��<ާF���0�\��B����@�Cl�kE<d�� ��]�s��;��i���T�V������גi�9�>{b�'��tF���k���r�׆U��	��EG��͗��g�$3r�|Vu�I��Yƶ(�ΰ���n)��l�`�Mv��ߙQw�;� ����[�'�g&R���uRP�����L�+�k�	k��n��t��6!�n������r����bأ����<
��=M
�Q�QNd#�⢆�1?S��;�MMXlxVHYEB     8eb     340R�O��7��K8���
�4�SĉR�����?M7��kZ]�+�F4�@�8�ͭ|�^=ږ��������aٕ�+��'>��jN���?{0=�L�Wn6����'��p(��]�Q�7ʶ�j�&M\<�]����K�������E(�S�3Ճ6m-���"pF��m�2Bş��2L��jfU~l����y�C8�<3�Q��
�����A�@g�G��M�h�K�@�l��r%Ǳ>W��Bzt�+��'ֽǸ|��b���S�B9
ى�7��M���=Fpʋ��y�}g�l
?��}��9$�o���f��4��6�n�]���@��!@r��_S��d���e.R�>�3�im�����>
"3eԗ��Z�h��D��+�A��FH��Ԕ��0 ��Qܺ
���t�ua�/��
,������>F��1V��/�{0�G_�"��C���_��Q����V~� �:����E<� o�⪘h�>�I����Ŏ�>7�D6� ER�y�}P=���$˃ ��K�W=�g~ 71�JÆ��T&�]u��G�l�>�3�<r��� �2��S��T[	�~���{�%ӜHj�L�;��e�T/־5ވs⎇��68�q�H��0�d��P}E����<;y��\�����ۆ'R�Y���V:���m%Ԇ���S�����Y�k�����cd7���3������k+W��Vƞ�D�֯W!� �E_u��IS�K��Y���u�Udo����	u�!�|8\�cr��c]\(3T��:��ia+��?j���¶��т�E,��k��v^T<�f�0�jfGr?��