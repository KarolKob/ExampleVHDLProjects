XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�7z���Hm��b�~��UA���������fEYg5t�ͦ�H������h��v+b���>��c�fw[���	, ���"Ƿ�����[��-����ܹ��}ZZ|YZ'i�d[{��f�������@d�Ь<{��c
֗Ԝ���X�h�vd��ց����eԯqH�lk�M��Dr���4;c��:y`�ө;���A����E��0�u�lE��Cdڝz�%�����lc�/u����^m-^�����U_čj���WZ*�Ȥ��ж�i[�?�p�[�D���;g�ED���ԍ^՝ %��6���37/��ws�V�ޔ�EIR���O;3�Ѓ�R�t�_�p�K	�w��3x�B$�|�;�Niy�"i��!��ϑ1kQK���$�ʭ	N���8����Q5[s�g�y_� �N��j�s1�[���3���[�w�B;1�^�u��"�5����=������rAW%�%����+1�SIw����.6؝Up\	F(=G�^����d�p�?��^�U�+إ��p�*Qr�����$GӐ����<^�}�s]h�����tއ�2y�!�T�Je�5	��)�6�pq8p"�),v���7`|���v�=yI��n�m�!�j��7f�=r�����L;� F�k1��������)Cy��|�v>�F ��I��!��c����b�����[Mu�Q�O�F{)�ԗX��5��8��l2�6�We`���5�Y�}�6^"�e���VM��sXlxVHYEB    1302     4e0F^��X��]芀�ȯ�lB3�J�8�!�P�K��}qn�n� ��4���͆���+J}榽�N��&�m��� UB�Fа�����w��h!UF�`U'n?9�ns��G��6_*ӎՐC;��jy����B��7��Jد��
�,\�R�< �R��L��C���u\�}NE��kЋiP�܈P��f�����J5+eV�����H�8���+�;l�/�uN�"y�V�Dp�@��U�0'�m��D�N���ъ�L�5yqv�%�X����<X�]�$uĘ��m6���:Nl��ڬ����t ��M�~~Z�vf��mrR32R.�����XsqH��EAf����E=yy�#��~?0�e��Ҁ���&��0�e�o���{%���M�I�������`4u����.҇�LQ	v�nr���+#x�Gѩ�P�?�uN�}����������}�H�EK1�G$L���\g�J��2:w��h`��Ŕۦ��0�/E�g��eܞ�ܫq��6�f?���<���jl�,����]�Y����t���Z�(Ԍ����q����$!w�)рȀ�G�]��$@��G���{_eo��
Q�DǙƺ?9�-p����J��l1gF�1`&ִ��7X�v|�d��ܙ�+���.������$}oK�*]�������y�<y�&!-&h���Lyo���Q�۱E����9��2�E&���'���Ti�����)�M���-��	+b�`��t��c�b��)�K/���C�����xt@�=���N�'�-�/X���.РS	[m^Z��Z�M��i5���V��k
����l�P�!*��y"���_*��D�Fּ|�zD����UԎ\��������9�8��<j�H��E��^�� "�L��]=�(��6�Q�G	�y�������-�:�crՁ(�Ru��5�*�J
q�{d:�{8[������܂$�Q�B�e
��4"��y*�Ƕ�9)��9��ft�0�l���jp*h*��kV2wЯD�ℎ@io�&y�7ܜ��/Y�N�w&��}�cưl�[7AIQ8Aq�����4e���:�1LRF�DU�j��H�}�Hrl��:3}I����҈e���Cp*�DGi|~�d
��vbN���خ��x�(�U�6ڲ�R����F��j�-Z���ȸ�"5!D9T���Z�AwX\�WC�.�;B�e�+�a�