XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9�7�M�Q<69'n�e`��ty��æ�X��G��eQ���)�q�$2��!$p��8t�!�]oq�X�2�f��$pwWR	�Py�f��bU.�D5�(�Za� uN1�؊w�hj�7 m�D��P�:�^!AH�b�%����y�m�,KI��ThOU��@���
��n���jLo�4�`�n��`�[{w��4L�e?����� �4A��F��w��t[�{ � 5
��X|��8f~�8�ۘ-�]�$���z����t��Z�6��|��'-LX�D�[! �����\(�HP��}bw�|`��r���$��0��WJ#5yΕ��;�r^��V���P$u��ݡ9��rj�hU?��1H#t���-A"�W�ⳟM�p�do�� V��$.i���h-G���c���X6���$H�}Qc[5�[�R�����so���^��Q�����5G���T@�A�v���R��y���_s�_H�"��Qb`�l6Ґ�M'pc�x��eo8�$
Η��oJ,����b����"�:��c�,g�b[�
��H�%b����@���U����tȉW���r�w�hk`�����al��.��Щ\[��vJޥ"�k���'����<S�1V�����#�����$V'\�i��d���gaTs'#������{�yel�Q菲�&xM�xT�Oc�nW@.��q����P�����Y�o�й�Nm�����5�!ۡ��]ue���^��Y���:�)ݸ4-@q�%����Z�XlxVHYEB    fa00    1960^���Kw��|U0P8g_�-��J��
S�z����-bf�h�C�/�y�G�u�na���뎖�q��(�8�Ŷ]	`��JoP�g��� �+��%���I[�I/�D��b(�8���7��pq����K�)�7�B�.Ls�y*�6�"�C��=I�W����ha�}�G�K��")6i����0��@�پ	�*D�=��"	1�e-�� �C��QN��$�'���'��"��K��qZ�i�&z4B�n&�_��{�,.nG4Y��4�l@F��z9��½��:�*�Ӳݻ��)��%GF�H��Kg�~��}�tM�F�9�]sL�=�X�yцH�!�����5�	8����Ű(|�h�Y�USP�t��+-h��*N�YʮfsO�X��;�]�-Ey�2T���"`� E��&im�����W�ಖ[;gQ�jK�8<gMs���ʳ�2�]X��l+�:��������レ�`]��^H5�d;�7�3��0$��,ل$�2\���NO� �����f��Ӿ|�rF��O��+�SX��`-�O��&)�"/f�Q��u�8�Gc���0�J2�����~�3I��4������n�"��2_J'�%3�g��n��|Z�9�Gav��,�fa�9?���57X�� ׋��*Fs�Y����c|xB�޹/��[���ͣ���)��A�G�����	�I�P�*d;N7���-�
w���F),��&�1��&��DO�g��S��i��oB�l���]F��D��A�bڿ��W̗��UD��"�89�pz<���%��ψ�p4?�0�7��ȼ���߸�詶���K�S��H�dk o��Y$(kQ!��j��r	p��Pj�*D�&�; ��V-��m���ִ��tҜb�a"�߭vY3�IQyt\|8����/�9�k�@����"L��SB3h�6J���R�֛s1,�E;��L�H�W��������	��MѬ'pѠ�*���u$�S}��C��^���ݶ���Oqq��]��b�_�tXg( �h8���J;s��h���t��Eg���Z>�c�N���s*o-7�%(�(-?s�C�f�U�N&�n�u�ު#��X�$�^�4%�'�噔�C�7�B����ׅ{Ix�I�,�B}7�䅬]��gV:�I��k�VՇN�w$cv���i/�Eh΢&��$�#�fT3�[���-k%Z�ek�K����a��������!N��t柠,�a70�)����~UJ�>b)ul�Xaݱ㙸��B�H�զ����C�si%꫒$%���֣ū5�uh'��,����W��+)(�����!%w���!�����%J�@��Ή�3UD,5hF��Ľ�d=�F���Ysɑ����ad�ae^ނ>����`�E�>I�L:Q�����2k�	����D�!L�k�]G�w�T��Cߡi�8I�C��q`�]�B5��4�U9�������D�څ�$'?L4�94�%�G�V)�:";"��L0Ǽ����Jn�2�CER����β�o:g�W����`�=�_�_�ٲz�qJ.�xLN����R��2���zr���<��a6�5�N �d[�L��u@���x��(���W,0"�*"a�a24U�r�e7b������S�HԠ��E@��X]�E����-?tc7��_��&�U莰�YW��;�yiQ�ʕ�zd��#� `��|���im:�acL'�5Ǥ.L	�=�K��p[7!���u��Ȩ�_�}���7���������O�\��&�U< 2��G��zYfbl6�hW�jT���;7���@���n�su���.�*{�1�+��/��Ź�7�YOr#�|W�����fD�)9�i��9K�y)C�������Q>�J>�fg�w3���7^��7��5|�����p�s��"�!H�m���f��HI4� �e���t�I�3xWv�0J���pef�&��9�r^=XBqK�wS�`�u�w�(#CM�DJ�`b�xg����+���tx�<ż'Ҿan��0�#��t�s�ypC��W�y���uMV��M��F���`͊��:u��s� �ڌR��$��[ٮo��t�cO�#: Fx ��g�c�v�)+��l���w}�vA���OC߂no��)���)�>��(¾�܀��da��f�_�	/��7i�""�[�7��s��3�}�p��c�.4�{H�䍟<E�I^�V�F5�܉��X��WT��0hO,ԁVS�[���՗Ȇ<l��>?ࡺ�l�u>�[���q�𑘧2���<(9IpzN��p�E"�$��YZ֨����t���h��R5ꗓ�JNW�`(�h3M�g���E�C;��Eʥ���v�&�Կr��Ѳ�� �1��@��t�j�QǗ(�D�U���5���|ʄ��`]M���;�,�<��O\(~d���!j�ToI����4�6�"�7���@��0	9�vK�Q��2l�	�O޺���c-��I�I�s��1���"���Wbnl�idmr����{��"?(����W�p�G��:Z���@^7kq֠��AH殺���RS_x
�n�MB�׺D90����0��d�2�v�]+������;�n�3�R�%�X�;)�)�h�u��-�A�TA>1�!B_�HE.CO�y$�3u��Gs:ч�s�)��)<��s����6*����n1��Θ+.�%	�����V���j�sβ���覢��NQ�x7�� u����u<ͫ��E�Y'%bE':]ݨk��C�Xcc4L�q$K�_�X���TB�Uq��p���w3�0��#њV������fƁ:C��~�֮;��?�h�΁2H��P������ax,��X9č\���M�{B�!�a��OWT��%.��v8��������������A���*A���PG�8;O�+�}�0��A���9�]J#��XCP�"f��Z>�\8�7�Lg��x(ʌ���?�	a;Lb�hFR�cx�DmDh`�N:�Ih��Y�p�+�����9ڑ�a�[��&'�g���w=�;�8+��5D�����޷�w�>sm���t��鳢0��[��[+7���DZT����=�dmE�
q��CJ$�i�>���~>�2�8͜H!F~Ð�YL8���ݛS��:q�N:��up��2"��Y��C)�WM����g� Wǀ�1�|�n#�3����8I�ŝ�P
�nB��v��g�5be��Ru�lV�7mFjV�����+nR^׍�;Sy�oC]>[�������v��l�BK�w'��ȽX�5q�<�8��NI[UH2����d�F��-�Y@��krW� !���S��2Ȼ6��MV�����ֲ��!w�*��'R��;��hAH)�����z|�Yp7Zm0	7¡��Fߐ��*��]��	F�RX,�P#E�P���&	)✘�f�uB���*RPF��0'ւYO��ؗ^�r��B��"���{о��T-��xөաG��=A�
��G��/u�RW[J�A�[ϲ���J�ܚIf�:��n�R�;L��\ɪ�U�t�]1�*�FT�-�E҈}9Wcf�$9�f�Ol<�:����Y">W��p���z��w�<�V~���� �3�Z�$K��2����53M��Ƭ<i]
��<�̼f�ט!�!2I�k�����qK����e�RJ��<�"�pؾ�FI�n�K��V�L�w���<4H�2GI2�f��De��K|��\��n6,����Q�U(.j(K��>���7b�EE�|�`�8JG@H��[U�o��_A����@�3�k�x����s?��k&�P��B�vfy�K
=[5�v�i񱿭��Z�+�?.7��oJ��G+ؤ��=)�j��h�H��5�L��$��lr�N^>�=��s�F��$�-�ė<T�USJ���b滪0$lU�$Ҝ�����c���#���wW^�P��h
s��������:����Wx��[yvfg���→or�t�J�#t:B��Z�Qڽg�%2G�/cz�FP�1����sR�L��z�RA�	�/u�1��	�Tg���ӝ��99+'PB�J"�	Fl;ȇ��5b�r�b���-��b����.3����N%c���s��f3��Cp�#����6cn����ʧ����&V<l��}��b�Ƴv[�����X��S����y�� ���.%����@�O$�|�p���T�'��$��Ǎڎ�t���Q�9������p�3@(�J��Sѽ'��a&,��X�},?i�v��:����v��ߝ��2G-���{݄*a��N�;��n�J?�䠮 �"y��4
����� ��ͭ��OGܖ������ս�~\�Ϧ�Q�Ʒ@��.���@��������M{8�&�m3=�t�(��͛� ŵ�"��x?}�g��������
��S�'d۲{��K��B|^�L��Ү�V���n�~.CRߊ(��rjh��	�8i���Wz�7��B�3����Z!Q�u�ZX|�4���O6�Wv����o�!�|��KD�z����'Up�E�%�Z�b�y��?��\#�
�ۏ���,4���53}�^M����m�L<m��R�,x�B��u�jq<��^I>v�ew{�a�����4���������͸vF�$_��D�����$�/.:#�Ǝ�v�N���џ��?<�i��-�ZZ�������-��NT��{^�H)��命-�8���D�G�dQ^C���}��F�::��'��r���a%�/�o<O'M\��z�yY��px�n��=ߞ�9��3��Vݻ��L;�nh����\K#��1��Yߕ�oRL\�t+(]�}T�%�3�A)�4�ESO��{/Q���x���E7��qwCpU2�]J{�E�{�k vn�Q7kUC�$A����Sª�n_Vu�����3ܥ�� �b
K�Dj���Hү{>����Og�*��B�� �&�o��ז�-o˳_BQM(��z°��V��6ķPl��n�����[0h�`}#�������ܻmu��MR�'U����ԛ{4�=Lv��De�-zH`�p��^�%Q
�ZQF��� w�}O�)�,�	;I��=��,=vI�J��^*6�,3+�g-���s���C�>����O11 ����
�>�0>b'��+�M�)�M�r���E?Ԟ>�I�K9��W`�c�}������E�϶*��Iq
1����#y�ƀ���9��2�Ɉ��V��?<�%��(��cz�3ha��?�W��k�|�v`O��Y>m�H���]�d!�V��(4�x^�v���"ʾJ��j|#���N6O�^s A��q��aVG�BI�-����8\7'��"I�&O%�\G�H=�YYYo�Khj�QA��,����4�A�1�T��ۖ ��|��#A$z�|���C�N�8���:�����M+�m��d����kފ<����c��ۺ�xs�9�U0���GW��;}��?%ϯf��&0���*Am �=���^��ST�'aO=�K2�RǤ϶d�2L���X���Ub�k�J�qW��e�	dL7�i�;J)+7��*|Lf�S[�Q�)]l���-M���$�������.4���"r���H�C�,4�ɤ����ROț�6�9�n�ïD��%i����V�0�4��3Z�����fF�}d�c?�U�ap�q������v�����'�I���<��k�lr9�:��Ī`0qT��|W�S�r{�m�f? ��Y3uƒ\�$q��.��¡rL�dɤ�Ͻ*��@p�!)�Oi0�R|l
�l;(��t�˦]���
�H|�]�B5s�D�j�D��ģ�3}菆�K�_�mW����b��Ixl�td�{�w,~H|=�7.�"G7���-��� ���L?A�%f�~l?��Ш��:�o��C�N]aQ�A�UB�g�s�c�J'�����־�E^�O�ԧ�������H۸�+2���ff���Z�G���T����o�h8�4x��!�;s�ǡ�� �5�趼��b���,�Y<�_c�>��P.!=5Ets�pw ��J�Ⱦ��U���6Ƞ���6#���S]	�J�7R#�r�/����g���9!U&�,1���<݂©�hq�AN���L��N#�5Z������O
f���FqV/Y͆�З5��@��G���rJ�=��b�������{>�]�V�����y+�o�N_��U�^|������??9p��T|2<��ZΝ��� ;��8c�/��(o�Q��s[��.(~����!f�A���>ɻ�@��>�TN�&+-Fl�F�Q<�
W�8�`�C����9��|��IVW�J���HỸ�!�VC���� ��#r;���]�}��f3���]�XlxVHYEB    fa00    15b0��$e�!󯬰 ū w͏fV���IK�Q���ǜ��
<��R�	����E�;�U�<+���x �r��[h�h���R�F��Ď@tt���ݵ���Xn
&ܤ������:?�Jv�V��,�")�CY
�Š����p��\Su��b���?�^��_�e�A�2����1T��,�kD�o9r='��<��P�x�Ӧ%�'�ru��r���x��m��Y#�JʮGv�vPs�Z�:n��e����d�r�nGf���l����-�g�P?C!���;�������H:�(X����?*E�TNQ�FZ���<�K�2��M��<H��^z��J���V%�<jFn�B��M���rWbRa┛��|�*���D�[���x�l^T�����O�E��E��U���o\���s7��N�{����ϠY=		��3	��y�5n��� M�
��եErkn����,�VWYެ%���e�[�L[�$7�+m0�d��t|yL:�ڑȶ��kNd�(�K ����
��qS�i�ٽqv�Ʒ`B�S+ rnl�<��W���xT�p��S�IQ�D�R7 l�I��q�Q�J�(�ۊ�z��1_0��E��E[��-�Y�,�g���(2���,���'���𕫆:9p��Q�Pح�{.U�K���U�{d3-�.��vk�E�=��v�e�^š1��o���ڛm��~����zڐJ������T��aٚ劈N�)�����F&��$�FDT^���	ڬ��A��(�g��䴪�'��r���Ż��0�??�E�Aүf���q����_#�|�����t�u�J���$�#��������ny����#D�:�#5��5�^2_�[
4�����<꧚�@��Z1ϗ8�혽�oa:Ȼ{�үJ��O�;�>�iE�����_�����ǋ�} �'� m߀��J�%{r�����8w ���� ����G*���������4�!� (�(V��=Iz.@����K�<�LҪpL�l�<���S��p�ZVpb��W��E�Ҁ���-?d�n}�v'"����d��{�M ��g�bCJ{n����2K"�f0)t�?�Ӆ���(��_3JYT�&�`�\���p�zM�� Fsi�ب��"��|�dEf���&���z�D���������p�O
����mW^��F跖`�e�X*�J���^��	^$��E(&��"J�[��Ʃ��%֍�6����Ť��	��Z1o{�8��xY
W�H�]���pn,���\>������5<�����6�+��F@�%*E������U��dC��̎���ι+�?�����-��=�����]�4�R}?S���.��ZG��N̒]t�V�:����4띳u��U��Bb"���M�.�TT`H��5I�xi6}K�c3���~�]���O�}�����|T��7�zZ->,����v�5w�qͶ���\���R�����>��0���	X���M�EqP[L��	��b�i�N��j��0�9#�A;�'��8U?P	�ꨰN�jƒ�OB��������tt�'�˽��
��U���!��/֬��[�,X����I��{�b���@,1�JQ�_&�G�w��a��ܡϚM�m�NF��s�v��<�t����X�x��y�ŏ���i����0�
���E6ḇ
�+�2����Ѥ�*��2�-�C>�����t���RM�qt>&^>"����jGѽ^�W��ſ�Voc�]_�|��ZJ�`_����} �]�,ǟ���R
z��~aA!K̏y���2Nh��W+�= trAP�^Pi��t�{˸�1�U�� )��7��5�2S��<$�cT�͈��U����N�(RE5*E�ߧ/�� ����}�5�=$íP��Z\53�9*`'�Á3�ݗA{�2��aƻ��N��iB�
{(J��]�aY�ÍG�'Ж�����*>7|/]L���O��mn�� N�`��t�ԺfӋ�틦����N�ް1�D �gK��w�8*}�#Y�|L�RoQ���R��܄G��P�7`�~���]I���*���m��(j����Y�
L��G\@�NBu��6�A5R;3��4VZ��>	�!�~�3�4�L;N����S�Sy|�fE��2��՚'F�!T;�,�� �o�B��nm�ρ}�YF�'D�y�b��"|/�`	�;iHi��o�vZ��#�H�$9iP[]�{��c*������-ni��\a �S�L�z&��!D�;R6nq+8J��q���dX3t�G䉯�dT�dކ	�����	�unTm�Ԭ����$+
�����������=�&g�P,<�'�J�L�XAyyҤ ���P���U� Wy7�Yk�)�?T��KXUV�Oe�r�j����^���}�1����E!�C��hB��+����ʙ�	c��*]6�Hs��R��`��>��%�NIR�n�p�G����9R2���y>hT:���Q�&D�Y~p=弰�6f3_m�O�A�!�ko|�����F�W �7�Ô��.��U����>���u��~�)�E�G�j8ݣ[�|���,�O��h��5_[+�L
�2M�������Q��\�^�?L���g������H��%Ѡ�UE����R�?X��S�!L]�e�Ջ��o�ff�T\=��K�����z��f��T��4K1�k�������p�֤�k�9�����#�X���
�5��̥Q����|e�	�/d[G��l�����Z�OȘBՉa�4h�i��`3�n^��Z*zz"���WR�����m6׼�]�"S�ͽ~c�f��Yt^-*�r�њ�I�^�O�ak�؜�h͏~�mR=����4�`��y�J�,p)ժR�u�<U�9	MP:�{=�S�H�A��Å��DB����qU6��>�0Y���侂�!V�ke��XC��������j���m8<�/��E�m�kZ4�g�5��f"�xFy���.'j�|�&��'6[l9.?����(ԕP��P�x��]���1@IJ�u��OHzuJy�G����٭Ա��v��\�U�۫�Ks�R��������0�������7���}�3)�qki�����`�)���O_6�:n��i�OL0����ՙi�2�׀J����6p�B��Z�r!6�e{����7������ש*��؝K.���:z��;�jH~�nqJ��}A��y�������Z�O(��ۏ�$75��l���iݢT���xЛZos�b�2�������~JQR��3�����:֬A�3d�nm��k�JͲ�6O��Ȱ�J�,��K��(��{&���Φ�D.a�x.�㛍+��Nź{"{4"��28�Pe��s�I/c{늬���w��&!���,r�ru0��g
�.����+��2��AtE3|��I	1���Y�o��_V��i�C}jQ��L9M�v@�� �ʉA��ൺ����@
 �\EKJz�v���@���SU��b��z�rI`|�Mj%7�p�'��s��������.�[O�PPQ�nb@4���sqc�
�m��4?_���g�qw�*��

=��s�	�������x���{�� �N��	��|�@vT�3crm.��VAF� �*�L�=�[�Տ�KǠ��&���)G�d$!�U<�(�n �ӂ�1�?�b��H�ߗN���!�(�t_%Dw��0�h8�����/�y M�����U��W^��.�+{�La�[�?+�����N&$.�ф��Mz*���eJ��e
�%%�`}�o���ֵ3Ė��_�6V��tf�fg�����*��<�����w���`_9jF��-�6JS��b�$m~/p��*�8FzL���ǻ�<)�@��Z����X~���,4��{� 戊?�m�u��l�W��ed����#��*�]\y(#��PA9�6����x���,j@�<H+t���v�k1gv�d��V4���fJ��6��٩a��¡�M�<���.�b��$�,���I���4�O[�0%*��� T��C	�`�%���2�s���4���sP���N¹r� �P�\�H~B��i�1�tbL&��3���ت��u�jX� ����Qy��O ��^B2R��Aj-���O{63���=F�<58��k��I�K��l?W;ߨK8{�7�0=AG�$��d_z�c~�s�"%�*A�e8<��v#��3!x�����LP�˟���bR	�X��7�,���O��`zd4���	��|~�^e�1ٷ���p���)��m��w�? �>���MS�ิ��A T��&�ٝ�0��6���ܘ�oa�2�c�*/|�z�E��_d�R�c|��c�L��S
����w��ڢ�T�SFHx��3˂m|7����e�u���"Z�9�H�����>�o+������{k�ᒝ��k�w󚐂_���f���X���,��(���M�0���$6^�<�{	��jvqyb�`��jp,<��O�0��2��@�W��cg��3G'��8M�C�GT��%!vz��
�S���&TZ�f��①���`&y���lO1ऌ@��qj�@��"<�Kb�q=�G��ʉ�C7��Yv���'4A���F=�;]a��� _F_̪��Ȇ�@��
�����& ����cݒ��l 8I�Cm���=0q��P��5g��[���mƚ���.���C9v>1%}f���c'1�8f��s�;㚘-���B�]���Ub46��uK���;�ԫp�25�<�QC�z�%x���+����%��J0*�%��l��xqt	���c�l-���#�U�g���Q�\��W|H.�yrix����=���Ё$�
��m{�A�L(��j�.~"��"*Oך��z3Ο���G=f6��|���4Zz�7O�6P�N���=���
嗫��xo���)>��m�.��1R}x��#����Mv2��u1a=�no��9��9�(R�hY���eClm�=ټ\*Oz��XF#�@O+p	U��r'���#�����B�K6H�C֋]t�y�y���{��"g5�n����@Wr9��6�J"�E����|U��|�$��ϔ�_Cb�*I���.yQ�	�}�T8���h{I} 5�j��!�Y���F>u���]޷.j�<2U�����i[�-?�	��y����^ �@�����Fȅ��l\��q�:�~v.)r�r�F��A�L��ݒ��|"�]�Sw�#$����g�������O�J��"0HI&g���a瞴o�|�����)�囥V�ϔ3���; �٘�@��=/$�O`�O��W�<�bԋM��^�m�g՘1��� �v�	�0��'kl �߹�`�]��L(��>.�n�=�1V#�^e�S�a�D�K�K�t��y� Ek�:Z�4|���{��Ȁ��-(�9d� "�����iȷ�XlxVHYEB    fa00    1600�!�y�cKl�C�yi�T�[�np�(6��2=���=Zޱ Z��=���N#kd�46���<��"th)��-��������9��p<gHk�F/���$���;�8¿8:��P��;�7F�M�ʼ�G������s�z�k��Yϊ�u"�  �W�\�Ƶ�ΰ�H�{�siH��Z� ��	�fs���ʉ��Q�U�pc��d�B^�3�&hܝs�ݿ�T��G�Mڐww�)�dM^����/]�y7HY��}��Uh��2H��Tv���}��$�CEI��cqVF�󭸴�\��f\�c���%:`�V;TB������M��=wĬ<{���R�RDw;�dQ6Qv�����v�J�:a�`$�[�#T�dHkFð�^��߶��T��r;�{�K���W��C���hMר����M��X�Ǆˁ���>�"D]ƣq�<f�co���*
V�NB;':�}��ʞ�޻F���f�|_�I|w�9Xdd��f�d�4S�$1iٹp��~m�Y=�ޅ�A&Q���������/M7WȪ���)�8��l����Tc,�SE��]P'�¼�����گ=��� ��u��
�f���6��Zܒ"*[L|�[�0RM!C�5�Y���:��5��da�/ ���!j����am��Oх�b;���`�k�i�Ԓ;�#��_0-5ܮ�J�E�`����w�zD�u����/wa@J��5|{C�X����R3��JK�����j��
������ۦO6��M��Y���2d:9! ���OfԲ�&��@9$�"�d�P�ʱ�F�3����k�����=Jgmh���������C���d�����M:&���O>�7�/�,��[�}D����_#��۴�,��{�,����� po�!�v�r�m3����Ω`�K�2r�R�~:h���燗c�a�TYQ�˗f���d��^i�!�f7u���ʲC���$#�E}���k��Y8>��P��86�0�o�8I-=+W
�]RP��Ă�9�j.��ʔ-+�2di��m����Q�Q>��/��?�A�Qnݼ�Nk>����PD�0Ζ-j��o�o��%;N+]0b�� <������6)q�e����W�d�l�pq^�tļ�O�31���&���BK{��6�'d_��4yd�[�m��g��K,�,P�Z��nW7$��w�jlꝦ%Z�tةu����+>�褞M��e���4u�V�W:��ŋ@��1�yC^�m��u���A�98d�C��Y286��¦Z�j�`�-/Z}t/�v/D�뜊"
�C���wrf<}�ny�����E�R7����8o�]~+͵�7����[{��0���{(�d5dA٠7��	������x�#�!��U�kExn�ƻ�rw+:-�,'L8�P���a��ܾ�����L��7ָ��NFaK�'�
�? ���l���/�A�n�gϖ&MWm/kWh�6��!��I^E�ɠ�o��[��s	%�.����$�M�G%��]�di�q��� L�(1�a#ݢ�8��ǲ�g`�ՁS\��<��ͼ�ɴ�B�>���$'��]5z�Hn@~��}d�5;���> ���$���P]�
'�8h_D�A�7��og�݇�7I������"S�?�}�������{��N���@*}Q�Nqɰ������N��ϐ
�$HM�ZC0�j6�u�!Q"ԠC+�$D��q��׬�n�H���3+���gZ��kA�A:Gmy@,�����̠�	Uί,����#n:MO1��[JP9�惨�x��MЗ�� M��+����$t\ڛ�}nұ��(ǋ�	����V?�WO�W�Һ��9��	ˆ�/���/3����D��I��8���Q�+�%�Ζ]12W0��ɽ/����!(�B�MFN/W#:�:9&v�洳�����h>*���[��Ɠ�xiV�+�N�Fb��bW�Z	+f ;/�f���2m���*���p���8w����>E��	�h"0]�4YqY�G��\|{�*���.�p�C�C)��`���g�GM̥T�Ws�J�`f\�ҝ	�]�J��lX\����R��S��|��D z�]xmF��,1_�n�}~�JY1F^q���%
a�e�Y��o}v��+�1*�4HV!l!�Ih"�|��r�2A�N�PVx_���{����G���b�K��.Px=)��76PUN^��Z�6 Y��9��._�iB\@���|��)r'�����]�,Y)(�V.͏B��Ɲ��B��96"�4�El[�On�&-fm��3����۬mC���A���JJr҃�EW�@�Lwzz��es_�]���3��[�x��G_���p�ĥ`-9	��U�L� �s�A�΅�$�.o�4
��	�Ts	���J�=D߱\*����i-�jƥ�5/�$(݆ �i�8�acb���ԉ��34\A`��3���؏�+��ɥ�h��Zm*�6��$�#���� �����e��{Yt��!��(�63��Q�/R�bqɜΠ+ �V�.�Ң��y�B@_�	��QQ����}�P��ı-b���)a�G=p��F?��R+�СL��+$�����K�ل�����(��	K��uW;�)�~J�(|���#Y[��Q�	��>�oܴ����)�J��VC~g�)��Wӌ*G۾3T�2�)P��o�����L��,Չ�"91[��1���Ҍm�L�=�\��t��QKȇ��+�[�а<}@Y[;�ׇ�Z�'D��3�	-cja����P̧�q�a8��.��4�?��>�	 ���

��KU�9b�g!}�wҴ�?�=8� ��mf\Dآ��7�~Ec'�NG_�¹��T��((U���N���t�~C�nm��K�󿘴����7�c�C���ʥ��΁�`|.�W�C6O̠zV�lE2̨(c[���вކ|j��v��(��s�CIxې��F�JzM23/�&������j4�ø|~P<p����r�&�=���*/���L;@����]X�����#)'���� c޺�Y07<h�@�CC���O�����ƌ���)"ͅ��/
�ܐ��Z��?��(9ȶg���X[�ē;u��)8���*梌Z���ʒ|���3�߉�3���ue��Z�S��D���{B��l�;���.2*���	����9$����U�89��B���%�ڔo#*q����Pΐ��5H�>1d��_�fTV�lQe/:��Sf��@5�}^���3מN�2�0�����'8]#"_sK�	F�]������c�@5�،�����*�Va�֥�N��{:.L�H?B�Q��.���.8�s^���6��M'q��S��0���Y��˂����zNo�`ĵaW�1A(�_�V@�s6Zy�{g���/D�/6�� ;�:&6ŷ�e~C�<�؟7��`19O�&�5�~�m�4��-�-r�����$J�=_���ZW�}��s�`�ԴSstI�!Yl�����E\�x�M�"yM�����YP��i3A���������-�0��ݰ����ڒ�D�ޔ*�u4�G�0��S���g���ˋ���|��t��7�nD�/��v��:;7�l���9'l�h�8_�C���Z`1(�Y�Ð�|���7K��f7	qIv�y��2[t�ol����ӽA14K�Ll"��g%�S��I�f�'@���䥍�|K�}�Y�Z�D�~slE]��"��q��%�k�L˷D,Ta�N�~�*A�`L��8-��iX�a��O
���<�8mr,����5�;��;�	�X�y�e�kE2��x�+)̀u�����YQ�y��Q��Ejv L2�2l���$ys�6�G�jR�����F�n��rrkv��S�
G����,�.
u(jw_�i�c���Vk%ev�]:5��S�)����)oo�6|$zD& Z�
уp�[�ed�+m	|-k�M[�fW��A��)�����X��u����7
�P�5��<��`I�$�|`�d�S�L�G�;��B��3F�f�/2�s"�� ��C���}{����6ϝcȞ�EQ� �O��<�}=P�v���I_݁V�ym�����K!XddW�]}�"ZdcRy8 `_�q�E-X\���3�&Ś|1��>:X|�<g�ZO���әGm���_�࿽�_Uh!L�<�W�׎{{�E�i���jK�w���Ux��J@ �����E�tn�}�h�� � &�p�#~��ɷ�2zH��jJܾs�*P ΒRvl����W� ��.6�:�/S��U	���σт��ˎ�{�~ �9�ܕ���&T� )ڟ�؞|l9�}u'�o�6�Xn��Yu{�GeB)m6� �<� �Wƛ�t�h��e?UY-7�kzJ�?a}�/b(G����!d�)cW�{y	��&w��Z��k�g0�
�~'���>3��ZT���Y����c���"0���Y�h9�h&o*�f0�FP���*��M�3GT�����ct��U�4n[�V(�|���L�S�P�1f�}�M�壟f�;���Z.ř�O��G�'�W~��Ҝ�>[�{�!���2�V��3=M��jI�&6�2ڄ�hUo���O�M��W(%�S��*��Њ$Y2�I:�t�.�ES�:��Z7V$����	R=M��~��OS��-�KO��m�����N]S�@P�	P���}
FL�D�7�V��n�'nҾ����S2kQH{r��G*����W�"�+���ݕuH��:�G,���XʖX��n�&��־ҫ~PkM8՘"��8����s�q��{�8�\��^�V�E�U/��>I��bL-�})]���)Ln���"fz�ւ�-�D0����0�	�4-KI���±�4r�Kj����F3A��C���{MC�D�9Q��B�ȫszj��݀��	��x=4�:�����Dc�vH�J�����bc���V��ḓ{�/3�B�6)�^3J�S#�R�!����� ��Tr�Z�%�m��W^�F��l��q&u�5��](Ir8�	C�M���u��̄�	�L�G{�X}��6�̣8����#X���254��>J zGa��3�0g��4���|�,%'�̠�3>�����̰��̔ �(�\�
=����.7�MP�$A�������5@2�puw��.���)����ֽw�JY)m�Rʿ�ݚ�Fri�eP�Oꁠ��USPǏy`'��Ż˭R�������F��c;6��J�4���0��L2j�w�]ݶ�YJT���u`n��s�PT������'!�\9��ݩ��G�nK>Q�����=*�q�>�E��rZ�B� ؤ|�VTl�"0�m���-i���w�ݐ���:1��k��1aX�H%����kc�$�H1�Z�Fc<�|��&�d�r@r	��X��~��9��29��>�*�7��g�����^8�|�k@�!��6�Ȝea��l��\v�0Վ<�U5���a5����v}��\�ӛ(Yf��Qcuiy�Ӹ��yT`��J����1�����<�tP�I�r
��\e���
3�2�|��_<b�(XlxVHYEB    fa00    1630�m��P,#��F<����w�e=_7�f�Q�Z�#����rof2�HcK!(}B��K�a�|����3��I�<1��ߑ����S��i���TJ�'�xX.1�����x�}�m����h�軸���`���J��ZG���_EQ}+^��R��a�m�^گ�R.�40 I!;C���i����|SK��ڰq�5RpFJ���D���K�>��uj���[�����`�����+�6�H�t�a�����6:����v�]莯�r�S��-X�dW�21A��5�|��$�;"Z͟���`�^0,�>�6�!�1V&bGE�^<���mmO��I�E����q�u��E�(��:���--{��\w{7�6���{�6�n�}�P��DCA�:���<͞�yKC�q�3?R�Y"�6��Bę�Q��$O@���r4��`٨O|8`zl� �ڮ�a�:3A���[yDԘ����>�2?`^�Jv���Ly2DkGKA\\�WQ�*�O��Ꮰ�ˌa��ўǓ��Y���3\� 6T%Hu��E�G:��`����7��� �D
�ia`5� A��d�E�֮ۯ�V����ƽhx/��mQ���٠~:hg�ʬ���*M{�?�w����m~I�So�b��c���>���ؔ��}L~����uJ�V�y�e��s�?�2��ݫ��GОV�>"O��#0eUcU�1�_9�QW��y'�Ӕ�. �߶� �
��q,?�O)[�;�p����1CiQ��Y��������.���������㿨I� ��fϽ��� ��NL4�a���V_c�Z����4^z/n�������٧8V�G����/�ɸʧ�u)�~�$WP^['������Zs�ԁ���%︾J��6l�o����_�`@����0�R�]Ai��t��/K� ��/��������L�����&^Qy�[�e�8�O�(g�q�=�����!\�
uږ���O���i�s��-�h/\焕1�$͛��z
d
ė�T[?L����T�4�Ɛ*�������_UP�Z��Q.ʶ�����V	�4w����2��m���!���ӏ:;�&GjP�r" A��y��M��+��0�fM��d����g�[a�8��6������KPG;�Q
�t�<�%����&��5�́4x��|I(�Y����
0ie�3�E����K>QBgEQ�od{��^�'x�p*�`����Iy��tֲ �~�-�@���=F��<vtD�V����V�M<�^���� Zh�5U9��_|4tO��x�0QԜi��	J�g�X ]�:20�x����Ҭ{�P�-�܀Gu)�'�%�4�Nst���k\H��x� t��S��1@OlE&��C�y�AɓRdb�3CO4����͑���s�� cg�6��D�n ,	�|��!r��8��9�??R��5�\�t����"G�h���	r0�Y��{!7E�d����(��W���RO"8Xy��̌D�@�v���k��6�O����D�
%��桹�qC*����h"�m��zV^�N�槈���P��r"9�����}�UD}��P^�]5bq����?u�4 �l������q�rS���>���\�T���Z�\y��F%/�M������^K^���UDz\���Pv���5	V�V�}3l��C�u��)#t�$�7���Eީ����<�ӸA}!��И_����Rt��TܤN�H�ySK�����t�X�L��)p^(HP-�;o��h�	�n�;8��fW���4�n@��t�b?3B�%�Q�������F��B�;;Xa��>z�@� <cV����{���f�f�����p�Q�@�B�O�DD8�P���?	R-�si.������_��"���L(�Q�e�u�C~eA�[SC����Ek��Y� +'��;�h@jogp�2C���v����^�s%��_��7i8`�����;��w�Y��T��i�+����e`eA��g5�ˡ�dY�0�<i19�G� �U�T��B��)�4k��|���3�ԑ0�C����v�1�^U�R�4������!X�u�f,�I�{ؖ�	q�Q�� ���(�H�c*?�2����ܽ�����xș��m�F}�����pl�N�$��̗8埀h�2�
�])�����TsP��N���X��%�U����j�B���|�A�WL.�HJ��Y�nvE���H���U��B-�F���:�� ��:���(�"����I��t�A��ShKh8b�g^ǣ�߅�Q�d� �-�;�Uى��C͟׹�x20۩�0��o�.���~x��XC�hj�g'�@�q�ƣ���X������k)ۂSS��/I��0�^t���A �Y?���+�I�A�h�/O��r�dh���K�S���n�7@���ߌx��rA��Q�^٬L7�T˾�*�?&�a[�G[���M-���x�g�d3:\Y, }��	��6tX���VX�J���?.�q�]=�EiQ���A3�	��v��OpU��͡]0([�� �)"���K��tmG�b�q��ց[6�dB� P��3|C���]���"���-��'�F��#�]n��<�!�}�*xY����l׉�Au�f��}HC6���w�B�����-;�ޖ}�`�p
$��s3m�(���-%"��V�hS�d�u�=�O^�H[�� �g6ˏ=�\Ԍ&#�{����v���ۘ!:�ƛ�eo�2 ��O5��K��)�B���c8�?�P���V$&�����ne�[�l�"��<>�v�c/�����c�e~;���$,t[Iq ��n�*R�7�&y���0[����5H����GH8C�5�YU
��X��_\��kz�_,�Z�Mk�ah��a�ּG���Tu��ڽ[�A����:�-w��s�
��ӛܟT���m% B�.��4s�,�y��[���e�r��B�ׄ��v3��.�?�@x��<�d��Npbi�0'=n�|��Ÿ=5(�Z��8���f�s�y��M���L4ρ�\ۑ{0;<�/hk����ݢS�i�W�'[)���b�����{�f���w�lRx��tS���]׵4��jzu�"k�ۄ�O{J��	hY��0RzM������f�e<���p̛�\$/T�h�k�����j�62����x��D�p_X�<�\��_N�>��?�m���ڈ@��|������A����H��Lk���x���:�@�`��̹)J�������ca�r ����::ɎJT���1��B�i�T�E_t�/�ZY'�7�]���Z�����F���\p�I�((�6�hTA���/���ʹ��a�{k�����l��_�3��J^1�".���e���}U���9�8�;f�*��00����f�?���k����m&��Ė�n���۾�ì����n��� �uFR�B���	?�.+���ND�Z�ڂ�������L�UƔ�-�K:����$lၣiMxx>
#'M�XP��L��l  |!*:"x�a���X�4���.�T��/������|�gpf�m�@1Y�o��G%0`����p���p�Q� ��\����O-��ľ����Mz��e�T��۴��=�7�(�\�8�����\%8GEH �/9��S7�{0��� ���,Q��\��+��n�QOH��:R*�q�m�|�0��:{��Dˁ'��ݴ��qAԚ��L&tᵮ�3��{�Z�;�#Q��VJ_�|�����N#�L�<z��h��U�K1�T�|�PL�(��"�Q� b�f}t���U^���{f�yE<�n&����X�����R�'���^W��{�K(�XV�ݚ�&�~7�)jx��m���a^݌� �_����<��V��}ò�<� 
�4f�K}�h���9��ӹ�7[by�+a�3H �3��`�s�����l2�D��N�q���Q4���X��(H�7�`�ՖSI8���V$���Y7���Z�L��}���>0/����Qm��}s�����Q{_�
��Rz�r����*��GQ�p����3�#��I��u������Q���<qb!.�X w>�΋<^現дgw�������K*	�̗��8mQ��]���KG�|���u�{⦾�U�F�o�z ���� r��KS�Ⱦ=�mp�2֩�h1��2�؄5nD�):�^d�>'��57����\�q��0p$�P.����Z#�$�k Ɉ���1�H���#��Py�X���Ӂ��o����z�)��ruF�l��w�� �kj݂l�<\p{Zf�v�Hfð��Hq������ڤ�|�C�Zi�mAx���0�>Y��ȈG��=R;�2�&�ۓ�� �޻]��6nd+�g#a�a�X�o1W����Q"骉t���:!�w�飁�� �.M!Aԧ����عz��m���w^�o��$)�~C�.CaJc��]/��Uy�sTG�}9a!��u��&´���H�^)*-G���:���&�.���-2̮�]\m�����e��&���:j�C�����̷�iŘ������5�� ?�C�F��W)�K�(��`��� I�I6�O��l*l�=��O^}ų�Y�X�gr��D��<�����;���+�-F9P�z ���xrB_���-�5 z�U�"�ϤΦ<��җ�T�8�}�Aw3�#;�3=�z@�q�[�����x�}h͎�MTh�s���y�*"��Pd�J�
1z���t�-Q�k�z��ޤZ��>��H�c�Z�����\_�p�s�`�F����O?�P��^��S!;����)#�R���쨝�½�/�������K"��̵�����Y�j&��ժ�Di;�����NbT�����ȷ&��K%�X���jhZ�VX���;�w��lf�X�_	���r��اg�#�������C�o�X��'M>��!�ڑ�y����цPv]���Ϫ�Ħ��&�\��:����L^i��5$��-�OE�N�]?��+�B�3z���fr��<�z��^a�@l�\�Y�X�a�gw)�=$��P�i ����y�8�D�{(�q�������<��߰9��J��wnlp�*9L�<F\}���%���0���NMa#bb�^�2��H���H6�|��h���۽��'��j~���U)����,��~(�.p��Z��_c�MC�I��®�3�?vSo;(�6��KDg+]�^��HoI�;�IA�aF�o�h#��p�&�s�^XoY�ڗ��Ѻ�/�f���5��;���m�(#k�����x�����|��.���?���B�ֻ�i��(P�^�o3z�X�&�v�b/P@X�T_0�Q��٬m)V^����9�?�!L9�C�D�@[a#����=�^��7�(!e��;2U����@�A8P�����0��F%ze�2���������J 	�w���S45��]�\�Ȱߏ��Z�+��������9�ɝ|���}���qU��O����tΠh�@�-u�R��4S���O��ݵ.��{��J�{����b�dq��l�_�R:E {'������&�XlxVHYEB    fa00    1620+�}�"���('>Ir���<O�4��=�j��M��/�$�|K��a���xF!�M7�ĕM6?}��pN+ø���/��ӣ��&A�g��K�vp�F��`.1L�Wܗ��s��V,A�^�\E��ݻ��P��{)2�5�:$@m ��hp6<T�t<JC9I��݋��Gf^*��#�����i-�V�^ǜWk&��{�� 8d�2Ef
s�7�|���x�Xɬ�<Q4�r�J�/�.��k��H�	qmO��n���~9�$R��.*�}��4Df��_;X^%��XBA�Il5i5m6�o`����/��)�Ua��.���$#�����(º6�%�9 Q$ ^�,� ��ɶB�$h�7ꑸN��V1ëȸ����Զ�_���3`>����� �Nר�Ӓ��U��m(*<QH�>&�;�m<&�Vo:m�[�_��)�Rtc�WV�py����.���D��.:#��ˣ�g̮����.���z�����]��9��0ebm:�v��<�|�Vs����J
$#��	YK�3x]>A��.�q5x��m�]�P^��X%&��=��2���O��mh�񠂓{w]�EU2Vd�nD���A�1�){��Y���$���>�t�4"|�)	� ����ܰ̊0`��\�~y���L�X~�A�ji�&�  ��!��e�TԹK�*�E��;"���c�*�Q�c���,��@��2p��%s=�ЧѶ����V��
vT"���ii�(�n)CCh�ůD�S!OB�Ə�V`���ϥ:���7�L�&(��K�A��;�웞�Ђ��f�.-ܿ�N�^_)���{+��ZL����2�=j�SI�{��t�-�yV {�a��s�;=b�u��'���Ke�5=��^�]��ӡE+iLsО�/�����|�Z��c�8zj�a*�'F*�jO�f�f�?�<��Pΰ����b����@O�]kE�Ht�`%��[^����G��@؜�� Q��a"C���W�c���r]"�@+'����9��9�	�SZ��g֊�U螣�����M�G-q�v�����IY�ǈ¡}D���$$@�����1��R�I ~�ѷ"�Ő� �T(��;�id�c���@=�c�֯b�9��c`�`���4�m�vZ���\�ޙ*�&P���41���P��x�u	�J�� v둑2�.@��z�Mޑ�nMzeј�ʎ�������$��bj;U;�H���^��³|p�E���+�'1��Kp��*�&]o�,h0dm���+��� k~�tC�?P|u_q�^��J��dȮܸqw>�-N�0~�y��f"�Ϲ�P$�r9h$�T~��0��in
���8�M*�K�5ó ��	�X�{,�"J48�����6��ř�|�C��x�p��)��G;�]�������;[1ma�&M/Z�z��6�PWD%&��� g�Ir��;�t.���S���K�j��70�1<Ϭx�h|��F��?R�u�q��Ѩg"�h�X�K�p|:x�=B�ն�����	qbv�w�`�4�!�_{^�DAA����������4ڳc@��|cQ��YtQ4�t��̟Or	�1��Ez?2��-����BW"!�𳲌�Z�&7�F)���*��o�$�K��!�R�)�3�$�r1��H�K���
òKuUY���l.M]��37�"tӉ�NA�p��'��HR-��T�m��o.��h_t�4e�=I�Xk�z����+��w�*���M�3�W��RZhy[��<��?�Y���ю��������G-�9�d���ϔ
�vx!��b�����*� �v?ȏ sF��Y���M؅��<�XI���H��S�p[��^�>g�ZJ~���0��Xq��?�|���	��mg��KE�� �k|�/�H���\sl��B�;�
"ʗ/|��v���F������u6w�إ~@�B7�7��� s��L/���hq�ĉ�Vc$C�"?Mc^qZ����͍��@8�	����pг=_Y�H��m	2�AO��������m�f����A/YF�4W�F����Y�j͸
��t_deɓq!��M�K�g�<v���0a	trp�ac�Q�M8�I������|�x�]D����mɚI6&=�:�T���e��� �;f�
E�"WŪ!	]��	��Nu.�ܾ\{I��+�����d
wH�/ 9���wZ���*;�����^� q�6"�bs�/M�+������o�c��(1N!٥�%Q����[>��Wۗ��%5]�U$�߰Qri���^��\6��A(|��h̴mS~T�+O��>�yaNNl�~�`��e�f@��gt\���1��t%H�vVYJ�u�Q��~,���@̏ i�@�$�ةr�u'I9N@BT���{Ƌ�y�M���qo��j�N�$���>���@.��F������4�,�;n���+|�������/q�����w�t�}�>�^r4]d �S�~7�4��gH���]��>��G:���TO��.���'`��#C�������ƨӠ+��+��v�m�M�w�M������}'	�	�^R��dQ��V1���+��o�YwBo=�k4��ߴO�����ϳ��K��F0{F��,��q�jri2��NL����A��ul,�"p+���[��o���N�_����8�x�� �}%�����4�|Mp�?>�ǜ�����Z�F~�%f�� -0
�C�s������~.nH4`7~�k^�㙗���,d�.�y��;�0{��Cu�����Oni�A��;(��<:vՐ�<��8�"���� ߑEh��/֥��W�OB mu�Rڥ�p7��Q�O�[K��5�E�>#���fᓑ&&]�
�E�܀����^T�z�:0�zT���Q�y�G��t\Ll�Q2ށ�
�2i�K��h<�D�xu���y�����jE��P�~��|�2������/T
��1��A��tZ`H���י{��˺H:��Ж�!�!:c�i��x:i�aZ��m^��M��4�ەQZ�抨U�?�w���?r5�iO�m�Yo_�yAVp��c"�?�6�vVk���
�k�0$ �cI����(�ɪ��ߏ�5��k�[_��KO5�3>�H�*��b� =9�J��C���M
��'���/Nm"�&m~<�0���2��|!��N�W�Bd��(&��oo	K���n�ǡ��ODᛰyD�@��@R��t�Wu��Rw9cO$[�|T�3�mD|���S*�>B��nmW�bd�Ö~]�:v_��j�� &G�^�[�������<�hͷ7)ɖ�����GBb����0^л��z3�j�:1�Q���x�z����5���cZ�=���ޭnE֊���?�}^�&��ayYr��_1ы��aA;��B�3��FR|Q'�q�(Q4�����9��5ЦQ��o��6�H(����+VQ	�n�[P5���I_&�8�����L�Q���KW�`$��ӚVt�̳p��<�e��`��'���хﮛ��c*���QI!�&�c(�n��g"�mk;&ۈ�-�;���i0�c�w����������m���4b���o�8(�p�}\��y�gL��:����3�f�g���RL��ɑ@�����t��ܒ3��Cbt�MN�$����T���M�+����L�=HePXӄ�U�7x��,|��Z���,j3ᡯ"�~{ulU_Vw..���u?��Ϣ�Y�?��=p��l(SMV6����2�ٮ�an�b��1na��T'[�7�������.24X^!��]9���ݣ�@�gGi�H�s3frz,��PC���DD�Y���fOj�T /3��ι�K�_,xߚEF�4�'8H*�wGZj&�H舻Kq	��
�)!�K��L��<�WE�o��|ߥ����2ђ��/:��Tq]L˿d�.3�⚧BU_j"��R�g~bE�0zN���xi@�fӄ�%� ����:J���'Xw��R�0���h�_�\���F��<.D�L�C�����ݯ����`Qĕ����MQ��m�t����Yi�)�,�}	3�g��vo���c�v_�y
��H�|��8�$��z���<�]�zP��sڱ�n�΂�$^jC��S�?B���(T�<��_˟5�ur��6��°]�?D��n��`)��7�U��#�(nQo��8f���1
f�o��vTH��]��r��%��y�����N-�:N^h�{tc��3�@��K���y=��礅��6�A����';�a�o�cs3�Z�F�u�M50�$�j��eP1=C��Ǒ�6��c�-�`�L翓�1��h�C3�%2����ڲ�����z��Y΁	|���_���/:�te�����@`������Ogm�C��dd_h,����a�}�����H���D"�~��#k��c��*�
��Cы�V�0���̑&����`��[��
�Rs�C�y?�j]�D�oD���^����K�4��������Ƙ�{�Fu]��^�ϻ��̐0��f� 1[��+D�F�-�R>k��!v��4e�o�/o�'���<>�P|k@�����5��fB�	��H����T�3�Kė8��s�[�|���ՙ@�D���a��gG(�˭Q�I @���chw�N��{>v�i
j�ԫ��y)� ��
�So�H���U=�6��e�l�0�T�l���~������h��{ɐ^��͡��0�եW�D���+���k�a��0�2�d-������@�m���ٔb<+UjU�,_1 $^���p��?5�^3�%�9�i�^�c?@�kso85�ǹ0p���5��zм������T$�g%GQ�9i��^e�U,����Ds��� ����h�P;���
8W*J��z[8�%Б�p�|�^A�% �w#�
O87�F��W�y�����T0և�fXh��'R�ᵿ�伻U�]�@Z�Y��$��iUq��h�>gFU.��l��Kdi������L���6@nC�[������?0�e�/�v��!2���iB	#��*;�/�v�s��O��f�3����GC{�2s���/��*�V���z�#,�j�;�6��]T�n�	��KC��Z�ld�٤ׁ����| ��cH�����$�ٯ*����hrm��!���z���z�C��m�����0��@�=�W���`�F�
i�t/�f�ܑ$N���,8��S�_�G?J�� � �{�1��Q��/��"���м��^!�����iW����4����X�_�8|�-!ӔQ�c6�]�}����!qz)�=��A�%��l��4�]� ��h:L���h�%�V��uLX��n��r_��,G�6��c9c7G�	�*��wݘ>�̃�> �Hx����Cl.���۶�Sj�� ŧ6�3Q-�Hi����RGs5�J�����nd1�܏2���	���W�m�£�`t��\Wd�H�4	4�z�u���[�r
Ko:�:w0�����&a�I���O,p�T�PXlxVHYEB    fa00    1630�h������f�d� Z���J�oD~9ծe�%�M���6E�xl�K:#�P1�J����7_v�U���4ͥ��05�>[��C�WQRҫ1�.���ۤ2�Ĺ���*4H�����=ٌ~�D�|u�v��U�=�����D��|����(QG|��ߐ���HH�n�6��)љ��V�߭�ն�c�'M�-��P�_���a�N֏��D���:�_4o ҥ�i s6v�	Q�B�Y/�s����X��Z�L�ν�o�4��
�v[;���-����(Ť�I��@�A/2�o؆z�l�y���#���a�N�3��;��˧0�H�}ߺ_on��Z�OK_��������
?�ю�\���Vvrh�I�����O�I�Zb�U�n�%%��c�婰N&�m!��Ds]z���F �(ڞЩV�RG���{x���A"-��>kb_/|dcC
)W�+:�t�
�q�I� ��~I)���#5�]�x��s�{V�i���m�E~_�
 ��X�P�5di>A��z���f�f����uA�E��H>��$����}7&�������EM��`>���I��<?;g��'W�����5Qlʴ#4��*R�|��`WK,V������Ԭ�4D��+WH��u��3�=���#�(��49�ty\)������o��+C����뙝 *���Qt�jUP�x��t��K���lg�Ɓ�7�-�Fy1.YF�#�X�ޓ����L!/2e�;�Љa�cݐM�Fm|C	���:Up��m��C�%�͖��9KE�n��ƾpY�U��߈�]U"F��'�u!v��j$��Զ��m���P>m��0��}Y�YR"Q%q;Y�Z1\��3���@tf)�n��n��,ގ��l��My�[ڈ�x*����F�S}��.twFҰ�_�eԺ������S0�a��9mp�Dۏ�}���MC��Lnw��<+�٢ԃ�C=�7rI95ס~�:����ti�:b������Wso=y���A�Iݎ�l] �-��
{עۦ�\�V���j�
���_��_�	gƧ�g������[����ڟg�_��T�&,��E<�$�y��Yh����mwi��\��|��@����F�z�W��'�x����ʨpqC҄g������Ի�W�qtK#?K?2'FiqG���BMSmsg,�Sߞ��>��\�Mu �e�n;Y��b�[*����M#��e6� L����ϥшu;��5��B���1���5	n�Mi5}�MFDj*�&-�a� �	�����&�j���ذ�9C�Y�1i3q���k��J��Q�(��9�=����\Q9���_���VY��bm��\;�J(�����(��<�#�	��
��������ӹ|��`'n��YG�=� ������e4����3�S����(/�}��,{ɞj��� ��ʍ������R�.g��u�%R ��[�ؼ����(�`^��bG�'ׂ���gg5�"NL�j�fd��E�AkÏ�RsR"��A��[6�+�6���Feþ?�O`򰈞o)!��D���9`'�"At��Pܚd4���v��g���{�N��I*���=�ҍ@�}Lp���W�9�n��p��W���-
�8��M��k# �d?�#¢wQ��M���ˤ��$�X���;�{*�����/\��p�M��WB�(�����z.@[���?_O�k����!`����li�iX�@�w�]����dLQ �ވ�W64D����/h˅�� O��^���~܇��A	q���������Mܻ�F�o���Wxn{"Xm�l��I丐4N��w�X:�u���s7>��it��x_�R	��	@����r�cz��ث��`��� �d���X�v�M*��%ؓ}ϸ�QQ��O����6�G�s�����l������O1S&�S�n��̿ADC��n���k_���ve�)[
�G�m������� ]��te��t�����we@(��֛H �+�^�L��M�T�+�ߑ��Q�SÍh�t-�0�{�GJ﫾��O<�k��	���e9A��̫2s)�
�m�xbd���Ђ�Z騒�p���~,2��?�֮��Y_v�?o8j�Ad�59�y$ִ�RT'�� �!���VyiD@�Vݫ�G/vw��[��l�#(7h��ᯩ5���=�0�œg�Z����|��Jn�Q1�)��݇f6��n�<>�S��gK^(�.�������<�=�^�1���3!�[���a���2� "2yXDn�0���@�p���]�H�!��	ON(�����)&����\"a	�5���䊠ʰ�e���%��*��1N���� 3��[�Ɖ�&4�e	Z�ᾮ�an� �G�(�"��M�T'7)�� #̨A�.�y�-�$D^�Ik�^l��\�U�g�uaQ�g�@566�#;/�O� ��Wb��aezI[6n��S�+q&X�XI�mwvBP�SwGÖr�o)����G{�I�Y��-��3|6Kݐ��Giʠ�ʖv�Gw]]ѫΠЯ�jԯ�9O�����{�:�� 6�'���L�Q�s��D��R@��}'��v*3"�x�o	�4.�g����I�|��i-�W�:�W���zx0�R��
�ā2�J��)�G����C��q�׮[;�����!�	�y��^<EY�kJ�͜��l�q�j�	�b��Rf��-�?�X�z�Y1L�{[b'�|������I��4������iP�� ��;���Y���}7UЄ�^z�&$��~Wb%::ݏ|�G�`{�D��S ������pb�D�\������t:���(]8�N ��m�Bn{+*�z�m�&��Eܵ��/G>��]����K������/QL��?�D��GF�Ǎ�#�
=M1u�ъ�!2��p���B��u��&0J_�D���	!���j��M����%�#@|��ʱ���#|���4�\�Ft�:�6�
^N��f�_��������h��<Pm���~��	�����!�mi��[^�#C�e!���Q�R�Uv;�S~�����80��ǖ{�9�N�bdi�^�q
S�:hJ
�4/�>ye{{<���Q�0W��Ɋ.D��侈�LU�z�"�YA��_{o�+ʲ��͜|֡�`/?�KA���)h^���s��$�1t����J~���1��(e7�2m ��G��K
N)�ر:�ؙ����֚�mm��8��u��1iY�Q���/"`n�woJD*�p�?۷��PVJ�e��cq?��t>U�0�6u�]�u�pl��.hC�r���W��P�@�W�ڍ��(�9�_��&��d	֏]��Q<���$�й�w��џ�B<�lc�Q���T�P�f�p�_�+x��&{�Վ0W��R$��9�U?�5�O��QD�j 4	�j��2cqc'U��U[���cW���T#*��jI����-�9;�f��r%�Ფ�J�&E��熌��f���\W�2<�p�u9C����֚��Jxiy35���k̛��`�@�}�3M$Kn�d�xL�E��Y�]�����gȥ��]s�%v���.M�]�g��o�p�`G��2+�e�\��Ŏb�W��c��@����v�m�M����T��;>\h�lB�`*/Y�ř��!��M�B@6�5�=����u���㱱>�f�S+��0h�)�r�߱Z��h���qI�M�**�π�b�nxܲ)ҵ"W��v�$�ؙ��F��[	Fni��$e�;��LYQv��t���Q���֋@��$���8=�\�sI(Љ
9Q�]$| R�������[BOѪ��y*ݥu0�-�.\9\x	�zA�omδ�[��F�ת��_��-6�H'5�j��������`���m2�@ ����C�GG���a$"���h�2�����EG�pU�^5ٺ��k��^n��"�/,i2�Wͺ����)6��������@)^N��'H�o�v��",z�d��l5v^��rtS��!M'��g%OwP�v��6t���.2d�˪5�V�["��v����t	���+�����z�)�G
���c���#zx��2���p6p��šVz�x�U5%E�YQ����j��yԍ��Pۡ�]�ȉUsS��lc4ICع����*.Z��'ۗ�_�3�ON��0Q52�	(�!�����L܃��u���4�] �Erb���ʕ���fil���Z����5Y�������Ρ��b]���Ft!�Og����M�a�qY�q��ZN�؀�V;I�뭷�~�>`�tJ��C~��:.�&'h3�W�u�l6��~m�S��g�5�x�B$gɅu���Ifs��i�L���ns�0d�Bֆm�經b#nsy��؝N�?&֎��!N�kgMQw���f�Jƈ���1���M����4�W�b6��!�͞.t~J�UNnU�'K�U��$P�q7
��K�.�&XL"�[\�����4<�VƦz�{���xK��!�.��⤻RP#�HT!k�{���1��>���aOr��Bn}B�|xM-Iu��tV�m���&��Ot�ҫ&��JaB�Z����u�o#I�ԉ`C��{�+�!3�4�4���(zU���;�h�}%���t	Ge����DCv
�j�ni�����,d׷��7E,M�@�Q�ph�Q�e5C�)���쁷��C鞝�L����7 j��[rV�s�a�Y�./vd�ZyU�e)�������^~�Ԟe�u	�>���'�8ѵ�1��
h�KM��WgB����4�uє��k����@
���p��d�!�p6�C���e�+��>p翼
�3G�#�Ȇ�$�cS|��v�9�x{���w	��^2(c��o,:�N���KN�۞�/>��U��LM�F�:8.}��Gi�\9�z��E����B������h���x����,�_S�|�Ry���5<��@��&�6��>���]�F�9*�;��Lؖ���]�(���3[���b��/�ŕ���H�{��۽_Es��ᝌ��<�������Ĩ݋�n�Z��ӀQT��)�YYS樱�#�$2�q@Q�k2r󈸿e��C�{�+Ւp�#��Q�?z���2$+��;�Y�����Y�H���mB�a�� O^��\���xK �Ebֲ���$_�IR�ɪ���[�3�)�O+��X�ߙZ�oM�.a�]n�Az�i�[�4�F: �KD"m�ª1%z���\�a�8jhi�h�m�����:�R.7_�4CYd�t6�J�ӡ�'S�/,0�H�	+����`�����>�e� ��`��oą$�P���7�`]{�����f�5g�Uq���$��ɣ0��&x8ƭ��$�˛e��Ͱ.�K�s(%�B9vs#Ԗ�*�(���w�R5�����]�#-������?;{�եl9�
�bwc#y��w+l�xƣ�UQ��U"�l��K�a�]�nTu-��@�j$� ܼ�öl�꾺�i���K�c9�&Qb��jS?D�+.���i�xd��붛�ᮾ~�O✴�H���X�n����~Y�;��0���v
O�.�O�J��ɷ�5�&�I�ɘ�*j_��AO�8��\r���5E
����)�*�(���M.�j���)=NXlxVHYEB    5a90     850-��ᦚ��l���^��J
_"Oʵ+i1����8me��z��l��E����bM�!zQj��pTN��5J�6�[{�tߏ<����ԷI[�VU�Q	���c=��gꁏ���tG��i|�Tκ��@��֌���3��p\H�S��%��N�<2ҕ��&!�^hj�cQ�ii�9�L�5���l]Sj�U�7��ݻ*ԗq��^�A�@O۱8��jԝ�r��;��K��o.��x�*I:k�(+�"�nSp�@�=B���s���]��;r�yLQ�hS��~eҌ���:ta���&R�d_�*Ξ�a`a��A�rOv�3s!l���3��A�@,��Tx;��$���v3����+Y�|�� ��cc-!t�j���3Cy�f�9ar��v�db\o�m�m<��7 �G���~�Bb����?y꫔�D6�X�+��A�Z`+]B��4ٰ�ò9l��a
�7�s�U���ibO�Y^��qﵜv�9� �6k�)2S�J5�s�C+jK�)��XW�Eh�w�d #�i	��XmM�҃���P��S%��&�3|�Z�W�Ïqr6jb�iz��<��|��ӇE0�%��5ܥ�U�����J����M��Z<��|h⣼M�}��l��A�d>r���*t�+�+L�k��f[�\Y�&��ֺA�8Y��vO�,��nI/C��a�{l;"[A�ȿN�=Q=�������lC}٪H�����rQڋ@z�t�$n�L?��l�C �{�q#�\��,����T	����O��a�ap��J^M����(�;�RPפv�/��h��|;k��[��!B��~(D7CE��l�����7�Tl#��!�闢_t�@�IaK��A�	%�0/�r'|�r˂���	����(��/S���k��8�3^����ƍ ��:�����Ԟ���ʮ�B�DT�j��ر�p��.��&*��1��EB"�}�jU�f�,� �\̑0�$�b2��0*��|F���Xi�D�����l]B���;�PI�[FV$����-��$��z�t#���{�ae/����gDK��aV078����}Z���|Q�!���7b�`�9<5n�'/88|��:6a5X��;�*��U�"���F�*%�]���Ei펗�E�5�����ڔ�4�&��C�P����l;�����E�&ajX���)�˕J�l�w������ ��#����]	�֪�~����Q}�).a3�zcui,g�x�/9�3 -�z���Ē3�qU79��lf V�IԊt���`mN���@0�P����hsy�� �U\�u_��A��mq����⩏���E&Q�쨛�9g�9v�`����^����ӧ��_�jF~�0V�a��
��3�F@��!���D���V#�;�s݈�� ��Ӏq��_v�
��Ͻ����븀����SV{���r{jNEft�B�44�k�`�=/q�S�i�[�� ܮ�Y�5p�������wE��Ek�45W����+����Of���:������N��d�i(��h�_Lz��/� ��s�S2�$`��c7P�rtX�"y��7��ƪ��n�����3=���Wy��	�C�K4]i����~%���﹵&�µ��ϐN��d�z�qZI�r�2��yW�'��6_��1fI��0Q����]x!3�d��3u��@B9��H��+xgy��O:�@��31 �o/J��~�wA�
@�j\+5Q�\5_����ė��7x�3l>g��� ��'�a2�?��z�cD�/�RR#H?�]��aG)���0�#��6�Zh��e�t�yŌaQ�D/�� mF��yes�B��;d,Òf�.u��Wa�5���AuFRYH	�iTE� 1�q0�B�{G��Ջ�`E �)����z= ���K=�l&�O�'�~&ة|9�($�bL:M�s����h���I&x��8�@���~7���פ��y_�Ğ�rkj����b��ƃ_�> B@�����d�[݊k�!Ft0mX[q� ͆-�$��ߐ��:c�©ꫭ~��oh�G�0@�;m�@�T��ٴ�@�uq�n�}Q�w1��M�~v����