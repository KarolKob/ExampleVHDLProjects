XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����?�+5$&I��7d8k�����P0����{
�w����=;ߊ�ϧ�%j+�O""0M�&�� p�w�$о�2\��DE���勵����0�RR��+bd�1��B�h�'r�{�l���V1�S���\m�O���SM���SpWuc���=��-�AL,����}���_�U�1�xf�N�C���ܝ�N���r�a�\����O>�Bo!`[�8�e�O����FPw��\ neS��>o�Y(�Z��Vaǚ}��&�e_�ٱlJ�n�[�l/�D~�\��s1��w_�o߀.�V��������U[��W-5T�u0�6��їK˙Y���}�3� q����?w;�_
����c·��l}ٲ$�6�+���QZ"Ե
-�1: �&�F�˛/퍗����܏�s�%�@C�.�v�,����f�R�����-It��3F�/��x�%�Y]{s$(x��`��Sq������T]�
�~��V�R�~��ȡ %<�@>�X6��@�N���v�ѽ?[�b�C�|+�t�l�7���W��źѹ�p��D�E�T[*�HYzM�0�Z��Y�c� �k%��=[��t�߲��2=X�e�Ϝ ��CGQ�[�W�������V�~H�[,Z^���*�:��Ԭ���	Ѫc ��z@��^�tyO�	��Y��u���o��K�g���律<���N'�'�hY0j�1�N��`�FA�����������Jl��&4�T��CTZ�8�"m	���|�%���XlxVHYEB     b24     3c0F���	{V�M�FJ�%�4��r�����i}�R�^yK�,���K���vMW~9h��ء��Y���l��m��`�e�j��,�bj,��+�O۴%C���ۥ��Y���wy�<fw*��m�z-	���l2�IX�.=��{���`�\Iʬ1EW�/�L�{r]�=���oDzg9�y7G�=�yF�q��ŷ�垦?�ꁗ�3�Uyh�s�ə2���#�@�'���f���欁�����=B�)��#ˠ�Đj+��Q)���X4�Ab����g���	;�����gxQ��i�_,��xY��K���
��O��Z�innQ��epZ�?���+iD̂d�-{j�v\��cO�h2�(0���F�B�� �,����rȟ����v�R5QDO���Jͻn�%��oia�M 󣠸I~f{Uʑ��f��u��mV�r\W�0�gF5�4/�b�3#x*�o�Xܣ�:/�ο$!��0�	I�zq@S�-zIs��r��SI:4�Z^���x�9H�k���d�8����ќc�N�����v����[.���շ����2bδwE)� 1F�W�W��O��(�#�)��v��O��(Kt�(�I�7Ѕ��:9=H!�dZ�c)!;]���}��
�M��ºE�s��8�[C�v�S�����/;_v\�0��E|W�tE�9�$�>H\Kk�Խ�w��ռJ+h>�I�J��>��.�%C(H�|D'ףM���� �$u�Uf6UT��?�c����nmO�M*���="�;N�3j�h6J'��*5HO��*�Ա%�e?ҸA|��#!I�p��+�?'�D��/�b���c�&\����G�
e=1��أ���u�\��];LL�@[�IA dZ�ue.ݐ���Y~W���d��p���5`�Ŏ!�$�LB?�ު7�v,\`qQ�W���-O�co(�z'�Z�3��i��g6�