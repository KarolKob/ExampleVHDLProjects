XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;Ԫ�Q؉CT������$~��Q#�9=�Y�Xmt���Z�`�i/�R� �dSxh���e󂿈>����9��"�6�?1a�z�uj/��^�ʷ�k����E�7Mm�1����·}6qx��'޶��	�N8sE��"P��(���&Zni�c��4�p�+�ƒo�Ў��"L��B��KVp7G~��/ֹI������bS���=De�x�Pn�A�kqZ����N۹0��X�|�:���
���h�Z�r��զ'ҵ {�pCym=2���\�6V;V�
�ћ�)��u"�o\<xjR��ˉ�e�H�� �K�9P��ds����ј5�lط���	�u8*&N�M%bާ�[J�V� %y����Fz�玀�֤bf�j��Fs��2^D�{�'5��G���l��k�x)-����uCu��kH:f`��|�-���_� F������߹���픏q�n:q��o���ZS�P)5��S�;�è�×�|qt�1S樎�=i���[��A�TQ[���a?9>� ����0[[���Y���[�~RP��ՠA6�>��<a�[��;<�	����ۼE�{����I	�2���#ѧ���������5Z��hM��#�"C�c ��?5io^����s�e�o�"�c��x����#[S��S�1��q=�C���yЩ�=񸥳@�뒱��1����Mi�02�g:Qճ���0���{���~�M49�[w����۔r��}�:<D%�¨A [�XlxVHYEB     7d5     300�C��*�êXT%�ߗ=���0;*Ղbk޵-�Q-��+'@�����>�/Į���W4��`��<�SJm�ſ�W�z;�issOd~�V��L�G#c>霜��kE3��g��:DjЁ3_��4w�B�J��W�/Ò
�,��5�F�>�`�O#��x@!ڰ�µnO�o�^�Pk���5i �7�Y1]Fg'fx�X���������0c5�	��_����v���\�ժ����d�\|�K�%���Y�|��E/g��F'h��-1���R�Ч��ݡ�T�Iڄ�,4�����=��I��H7oC�x�G:9�}�?z{>$/x�Cv�"�,+��{����\b�a,R��2�N�X�����V��z�Cs�~NaL� `�"|jp;=�;�$A�� ��b9�u��v$
�]��^�6�������2�'Y@�Fp:w������G��� ���en���=?��4Gv��+���&Utlo����`
����%�/}Ә`"�0�-��e��ckW&��W�Irm�Y��cGv�gb�c��iq�=��j�tX��ʎ-�u�yc��:(��Z.WI�?|��a�&�vƜ,�;OA���	���pu�rd}۝�b�����q��f#8-��ߋ�� �]¢Z��o��3���d R�I�/J���PQyf%bd#{��{Xpˎ��h��P�{)���nT̮��7%;�4^�&l9�U0��P
� ����,rྃ��8��
硡t