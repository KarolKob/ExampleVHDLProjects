XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P���
�f�}1���#�w(��2e�o��9F��.�k9�z6��� �s�|d������7���W���6'�l��h�E�E��hc��*�q7w.�Ao�mx�V�u�Z��J�R:��ў���py���lxg�qق�+�K���(�x��m*  ����e,Oh��k�PV���1� ����M�=����W����Fŷ]�Y��<C@�t.�2�.�ǘ�s,����4ۺ�E�$j��nN9��.^�#�<0�ڀ[�J�mtc�$9��� (��G^*���91�ʩX_}c�2�C�4R�%F�I�������p��al�:v�/��%!��l��^�@����d�	�9�ɑ+����I��p�����.F2����/�h�o�؀(�#�0PN��������xV��e�xl����/�p��1���Ğj�d1)�]��\�߽�7!�� �pu��t�����.��/�;MO<�}���$��f���s&w ���D�>�ՃW)c��yO ���o���R����r2<��u��>��pp6�O܌���{�P�`aC�3�CZ�,�ؕ�BU��kǏ�6��#鿳�r��ۅB���B�������Ȃ`%&��C)on�<�������
k�����R6�Yhjfy&����,�*}���"mx��������)�J�d��:�1�Tڣ�SoZ,��t%�}�1���m��ʅ?��a�,ј�Q9f*����n����#T���%9��G<���PXlxVHYEB    b892    1b20�߃.���(P�o�Oz
�e0L-�3��=��t��ד��4��x�Ujt �R���k.�I���S�������QV���eŏA5_��\����jL�%����5Ќ ��=p8:6?�+��$=?���; |�zR̛�-�}���=�U���H� �O�����b�*��q2(�m��(4e�6�&"v$����?�O��[��"rj��|��?�*7&o���ه���	�r����=r���Ʀq����)(�6i��6C+���~������+{g�5f+<�\�^]��@�TcB���������Sbg;��1JC7�v�%��B�ڬކ�����کCu�k�w��-Qr��+� X����·ܑ�M4��q��FR��A�="��N{�{W���vQ����N��G(�݆\XrMQ,~����G�nz�l(_������u�!j�3�>x3k�EC�)~����#���x�r�S�Z�KYS�Ft5 �����1Ts�$�5��/�P�B�8[S0�$��ˍe�¼��%뜮ȭ*��y�Q+���N�03�x҄ck���i�
e���p
�vij���G�x�������]��K��)�?��'�%�R�M���稿,��GߨD����������p�=z�Ȝ=l��\򣆫�����M-=�i�����)��ږ^�f�uJ�qT�Ym/�OJ�uϟŲ �ì+�t�NӬH��=�7脇��� �~j_,�}d���|����J��$���%Û�0ȍM�|�v�_�%����Kl6��S��=�E�|�1��Y2�{,�g�[5�x��wе:$G�d�M�J��s�r���O���:`3�|�8�y��ۘjZYƿa�C��`�'��!w���?�2N�GU��Vj�X�����dG�_�Fyg$jz%�����_<� 1D�̴m�QZJ{+���S|�!,?v��L�=ily�m3Sm!4e��=C�̏!�PƄ��G�Ђ��n����pD]�t�$~V~ux&)L*J^��4��ƌ�9���`k̘V�M�|���Tį蟣�p�[�M� ߄�L�gJ�N�@]Y�R����C�2[�"���J�ȡO��[��[��6Є�b��|�V�Q�Qdʕ"��y�������䮄�]�P�/��!i{�3vE�ja�eM�ǲ������>E���5F�B(u�$i����Ŭ��|��w�:�8�ɮ�
��@���QŃK�8֨{��8��+�:y�|���G1�t	�S�V��>;.���|/�H�ȅ,�s�b���K�j	��<>'>g��2@`r��RvD�f��{?z~<yV����o#�E�S-�����W��;�U¸�T�l�bh.M �8�}HR���0)y2O��	z��qᾝJ�a#x���1��i�h�ýeS�x�?��1[.-*�R��J@�ʫ�B+�7����pKV�[�hA�e%h Li����S�?LNڴg���ci-���t4����N�*���;f�9A�¶����֠�k_0��t�zQg`�}�3�J�2���\����.�`gO7����ʒL�X7q��=�wS�4��F ij,?0�����Fc#KR�r�JM�~oY.��nV� �P}��&x���� ���,˾
�� `'@+PV�?@v�/��}�Ͼ���7����7���RR9����-F�Qk�5���[˔��>�(w���ߖC��O�+��P�nL7����]ur6G��HP���`����wt�Sw\����ے�=A6��&�1��3��O�z����ejE�t�Qr������zko4�-�;4��?��[2>�����z�|�)83K=1��a�q��R��L�R�W����M�E�&)]l0��=�DKO�C�& �@�VSE���y&������^����:̺Nސ)蝐b�U|��VQW�L��P�.�_�6�����ϥIlf@�B�&*r�V���}��=��	^���S�ĥα�@�,�m��L�>�2#���ha�Gu�F����t�a9	���S}�����{Rby�sh	����e'�Wd2A��g�{|��=~�G���o����WCZ�w-z���������k+2�/�D>3 ���L�pK�>~��R���1�F[��
�lù��y�i�ե !���@Y.�W��z��gH�?[�xiz��;�y��A.FT�����/�v���b'������$�Hٝ��QGp5b��!��h����}e�`��w�*�l��}���
K�Z�WٺߩO�8s#�.�J���Wذ���^�W�01p�E;4���=.�D�\��˵L�N��g8g�y|�/֦���brϚ���7bXn7��8%����>�p�2u~�q������-���"�m��PkA��A&#��	ygG%:59�K�9_Xg��3�7.85�� �fa1%H�˶��^��f�w���S��ؓӥ(���UdN(0o��#���:���xO���}0}���CkI��d0<��+�A��f����&K6fH���B��X�
�S���\����A�;���,���]��4��))d��S?���������Wpgϫ]8�>�Bw}Db�̱��B���◛a�YЈ�J��W��#�*�ư^�����MF�h��ٻW�LhLX�F��82dB�U�qk�U%c��_����J~PeY�$�$ʪ����N19�F���햠� �i(,m��}<���2��4Su��<-����ji�h���7Ӣۨ���Cb�{<a��~�w#����&`���D�]Z�Eɼ ��^�U~�ަ�����g��l�l?Qpջ���G@�~�83�3)��ݢ��HL~�j�{���՚������9���q�p5q}M3H>�W#����u)��aRu4f�1��������K�v
>�Vg�d�ڶ�����gLx͘7%]3��>|8�B����~�</.ٜI?_wT��Dɼ,E1���g�;ԵtJ���I�.D�g4�V�k���=H����`ؽN&�NA�J���{7�x6�7׉�|�q������)�[�j`��j�k\�bM	s��Ȕ��F۫�u�{�d�[{e��o;LX��K5�9��.&d=������������y 8���
g���eDuF`Y��s���4��x3eN�a*����2������|��9��:f�5?i��_D�hׄe�Q��G���ķ/
�B�eo�x�������i��м!
0x��ڦi�����[Y`�ԱP�B1%�������1|���߃K��J��+o�=�<1z�U���iK7�4�Љ��e;&(���$b���8�Cv3 ?#�W~WE!7���6}��������)tĤ�p	���<ɩ*���-�YPnJR���}��e\R�M��;�\��4;`t�H�Z}J������̒R��-&K������AH�����Prn>�"��#*k�7��Q���ƶ�T-����o�A�oϐ�äVn${,���-����������a���3˾���-��*<W%�|����w�����M�1H	k\nH54'n���p�	��~���T���.A1%n��-��;��&#,;Gj���P��L����\���+�A�)�}��$N����-N�0�Yp��N偉��_z�'yXU:ϣ2����Z0��֪!�,�F���͸-[b�%e�4�Y��ؕ{��2�1����J�f�D�Øf�0��h
'�F=�b�=�p�7ӄ�fٲ�Z3����Ŗ���١<^�E��0������έ�UpjsZ������}����b%6T.[m���9�{׶��ly6���At(����@�5�+s��\��ϬR�3��6q��|����~8k��ĘS�E���v8/��D���hK�i=2!�sٌ͋���7P��Bt��?)J��Gl�Ϸf#�Vf��GJ�����G�8nV�wz�ڕ��۟�_6D0���#Hȱ`�q:��c��cax�z���\�����t/�����_����_1��&��$RUUT���S�&���dCי~��A@�ɣd��y�������x����x�����*�D|k��$�s�+d��d��t��AD>^��U�w#�,�n�'!H�C�!Z�(����m�AbP�?^��] ��%�7~�/�� ��B�K�*�*�\b�>���e�M����r�L6���C��}?�	m޶n��|2�u�u��2kC��Ӕآ�;	$��|:1����T���?6�����RY��)�$6�S�s�Ώ��%�]vҎ�|��;>��D�� ׹��5J�U^�� K
Ž���~K�P����!(L=w��q]7-7|�'��bSl XEY�T��qQ�IĩІ��,�^�o[�p���9(o�Z�
ԵT�F�	ڡd� �0�����W�^���VZ��PL���n3�Qy-��AQ���)��7�����y�m���>��S�O0���35
�r�V�^�Vsw��Y�O��J¹ѩ��Wݫ_8U��
KM�@VZ��� KӀ0C8�L�UI
�����;�3fe��!�JP>n|��d,����Ɗ����ق^��ᰙ�~ptM5�@�w6���X�IQ��{���Wz�T��,T��a������v��P3j�B#��`�oA"O
WD�� ��n������*4T������u��$c�L�X�t�]!A�*V7�&f�?PI�/0�J:ƴ�ŗ�G�(�sjA%��3�� ·�K\�`O������ 2�ef����>J�2^r�9DȿY΍q6���e*<&s�O�,�뿢��K@����la����e�P=����z��=g-9���Q�C+�u[�� 5��aUa�����n�3���*���g��v�zGJT���f�]��j���VX0�����*G����W��`_RE��F�`�*���O�J(�]�M3�Q�O|�h>�aS��@�ƣJ�����b�a����'��+����ʵ�0�S��ZT\ߞ�%W3̣�y��V�'A���I�e�P����6�5�����G${h���γ�w��p�&��S��\֘�<���À��oh��4��c��"
qk�YMZ�H���Q��UD�R�F���~_B[`O�9$��J<�'o�.g����ۤ��i�bL)M���GW�&-��u�BReM��.�!�#K���cՁo`ݨ��E�K�_0�UU��z�d{�\%X�H���,B�K��2 H�{N��	�W�-�y�B��K����E�bu*�ptI,sս��ޜ>�>:;�P0�B�Ϸ��f��E�B=���w�������!���l�!�҅Tm �d)�� �?+#Q�'eRo[���=�:��Y��*�L=���F�v�����h�ĕ~�.��d 	���L� [=�~��na�W����,�MGT#}�;�E���(-*���&�=��Ja֤�Xg%g�+o�+UK{7���p�`)�<Ӆn��H7;Ϸϣ[t������Y�4,��0g_�f�2������jU���ؔ�]lOɛ�E�h��3HJ�?0%��	ښץ�W!�g��e�B��2c70��F8`#��z��Lo:y��3o�S+B~(�=5� �H�x���B�!;xӂ}ou��c=���*{T.�b,�[��G��aQ�P� �>�6�,_j�"~��	W2."V��d�I��Y������I4�DE?.�!�r����b��p�u���VI���ف��&��;]h���Pm{E���
��%\R�諰TI�q���w�S~s�Rf��sj�ͣ'q^q]j���}��IT�!R�tS���8�tu�Y#�����6���l�uQG� W��O��3Μ����߸�~�� (1��e mX�+�f��1q�!�-��@��!ƨq��7m0|�R
(��g*�" ��W,�Vgm��Ye1#3<�L?���Ny�u�?i��NC_ժz��h���x���K��$	���Lx����N���7�4%�P�ǁ�hb����?�X$�?#�,�X-?�v��\�ǆ��I�`'V�H95����i>�o�L�sd�	��]��� �QA>C*�,��x�@Q6Q���'#ҫ���(��=B"�~��d�$�ӽU6{��V��7��'���)��'�@#E5��'���:h�>�M;r�
�@�����RE���p�Qa����xoS�z*���hZ�a�>�K�����m9�W}< ���LI|Z�y��Dů?
=�c7\�p�Ez�E۹.$�%��<ު�N�1��S�QN?�QB�m������l� p��cK�W(�	�����o�tw��,��;"��� ft���8 �B�R7�|r�8o��Ͷp����������W���鈈�� ��h���9�ڗ�!n=.��� �`0p7��GɌ-p����0�ɨb���c�@S� �jO@�`P��n��)G�b�1��j��*/�E�P�F�a(����5k��U�qv�sb.�/�`E�qa��]�X$�ћ���T���݄T
�����.d������fe���8��9��ϣ&wk����{����2��
�K�@j�	Z&�:�š3Z%ma_�GG��b�"ɮ!�d_H�@� �S�A�0 �=���x�n��}E�ԃ4�hʗ �(q��j-�=�[��֋�(����*}i�b��g��3�d�8ٞX����
B��3�MD�퀪��B�q.\��N!��ES�
s�1N��=�Z���W�#�����ʾ�����	��l[���aڳ?�S�-"�O��שǶ��H���x�]��Wf_���v!�)0л �V���]�G	�3n����[@��؀|�e$�#��